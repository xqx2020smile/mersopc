module mem_rom_weight_out_02 (clock, address, q) ;
parameter DATA_WIDTH =  32;
input clock;
input [9:0] address;
output [DATA_WIDTH-1:0] q;
reg    [DATA_WIDTH-1:0] q;
always@(posedge clock) begin 
    case(address)
        0: q <= 32'b00111110000110001001011001111011 ;
        1: q <= 32'b00111110010110101011001010110100 ;
        2: q <= 32'b10111110000100010000110100111101 ;
        3: q <= 32'b00111110010100101110110100001101 ;
        4: q <= 32'b00111110011101101100101010000010 ;
        5: q <= 32'b00111110100111011000001001000010 ;
        6: q <= 32'b10111110100101110000001001011100 ;
        7: q <= 32'b10111110100011101000101000010010 ;
        8: q <= 32'b00111110110010100110011111110111 ;
        9: q <= 32'b00111110011011101111000011000110 ;
        10: q <= 32'b00111110010000000101100100001100 ;
        11: q <= 32'b10111101101001010001100010100001 ;
        12: q <= 32'b00111101101001001100110110100010 ;
        13: q <= 32'b10111110010101011100101010110100 ;
        14: q <= 32'b00111110100110111000111010011100 ;
        15: q <= 32'b00111101101101011011010111111001 ;
        16: q <= 32'b10111111011101011000101110010001 ;
        17: q <= 32'b00111110101010011001101101001011 ;
        18: q <= 32'b00111110111001111010100101101110 ;
        19: q <= 32'b00111111100000110010111111100110 ;
        20: q <= 32'b00111110010111111010011110101000 ;
        21: q <= 32'b10111111001000111100010000100101 ;
        22: q <= 32'b00111111000111101100011000100110 ;
        23: q <= 32'b00111110101001101110010011101101 ;
        24: q <= 32'b00111101101111111111111011101010 ;
        25: q <= 32'b10111110000110010101000111110010 ;
        26: q <= 32'b10111110101010000110100110101111 ;
        27: q <= 32'b00111110100101010001011100100111 ;
        28: q <= 32'b00111110100110001011110110010001 ;
        29: q <= 32'b10111110000010110110111111001011 ;
        30: q <= 32'b00111101110001010110110000010000 ;
        31: q <= 32'b00111101111010001101000110101101 ;
        32: q <= 32'b10111100111010010110101110100101 ;
        33: q <= 32'b10111110010010001001100101000110 ;
        34: q <= 32'b10111101111111010001010011111011 ;
        35: q <= 32'b10111101111101001110010111101001 ;
        36: q <= 32'b00111110000111011001000010100011 ;
        37: q <= 32'b00111110000010011010010000000001 ;
        38: q <= 32'b10111101111101100001100010010111 ;
        39: q <= 32'b00111111000001010001100111100111 ;
        40: q <= 32'b10111101101011011111011111111111 ;
        41: q <= 32'b10111101110101011001110111010110 ;
        42: q <= 32'b00111101101101000010111011010100 ;
        43: q <= 32'b00111110110001001100010111001100 ;
        44: q <= 32'b00111110110000010001010101011111 ;
        45: q <= 32'b10111111010010110011110100111000 ;
        46: q <= 32'b10111100101011110011001011100110 ;
        47: q <= 32'b10111101101110001010001110000010 ;
        48: q <= 32'b00111110010111010011011111011001 ;
        49: q <= 32'b00111101101000010011001111101111 ;
        50: q <= 32'b10111101011010110111001010100000 ;
        51: q <= 32'b10111101001101101010100111110000 ;
        52: q <= 32'b00111111000010010010010000101101 ;
        53: q <= 32'b00111110000011011111110010010000 ;
        54: q <= 32'b10111101100100011010000000011000 ;
        55: q <= 32'b00111101011010100111110000001101 ;
        56: q <= 32'b10111101100100000101011011110101 ;
        57: q <= 32'b10111101111100101110100010010000 ;
        58: q <= 32'b00111110101011001000010101010011 ;
        59: q <= 32'b10111110011000101010000110010011 ;
        60: q <= 32'b00000000000000000000000000000000 ;
        61: q <= 32'b00000000000000000000000000000000 ;
        62: q <= 32'b00000000000000000000000000000000 ;
        63: q <= 32'b00000000000000000000000000000000 ;
        64: q <= 32'b00111110010111011000001010110100 ;
        65: q <= 32'b00111101010101000111011100010111 ;
        66: q <= 32'b10111101000011100100100001011110 ;
        67: q <= 32'b00111110000101000011010111000010 ;
        68: q <= 32'b00111111100101001010011101000000 ;
        69: q <= 32'b10111111000101000010010011001100 ;
        70: q <= 32'b10111110010101100101000011111110 ;
        71: q <= 32'b10111110100101010010101111011101 ;
        72: q <= 32'b10111110100111000110100000100001 ;
        73: q <= 32'b00111101101010001010101110010100 ;
        74: q <= 32'b00111110100111000010101011101011 ;
        75: q <= 32'b00111101110000111010001001110100 ;
        76: q <= 32'b00111110001011011110111000001011 ;
        77: q <= 32'b10111110011100011011011000110101 ;
        78: q <= 32'b00111110100110111001110010101001 ;
        79: q <= 32'b00111101011101100110100110011110 ;
        80: q <= 32'b10111110001001110000000100001110 ;
        81: q <= 32'b00111110110101111100101010111111 ;
        82: q <= 32'b00111110100000001001100100111010 ;
        83: q <= 32'b00111101101001000110100001100111 ;
        84: q <= 32'b10111101110110001001010010101111 ;
        85: q <= 32'b10111101101011010111010111000010 ;
        86: q <= 32'b10111110100110000011011100000101 ;
        87: q <= 32'b00111101100110110001110000101000 ;
        88: q <= 32'b00111101110000011101101111010010 ;
        89: q <= 32'b10111101100100101111011011101001 ;
        90: q <= 32'b10111110111110011011001100110001 ;
        91: q <= 32'b00111110011111010000000001101111 ;
        92: q <= 32'b00111110100000000101111100111010 ;
        93: q <= 32'b10111110011101000111100100101110 ;
        94: q <= 32'b00111101100110110111100100100110 ;
        95: q <= 32'b10111111001000100101101110001110 ;
        96: q <= 32'b10111110000000000110110010110111 ;
        97: q <= 32'b00111100100000111100000011010101 ;
        98: q <= 32'b10111101100100110111001011101111 ;
        99: q <= 32'b00111111000100111011001001110111 ;
        100: q <= 32'b00111101111100011011001101110101 ;
        101: q <= 32'b00111110100010011101111111101101 ;
        102: q <= 32'b10111111100010000100000000011101 ;
        103: q <= 32'b00111110101100110010011110101001 ;
        104: q <= 32'b10111110100010001000011000100110 ;
        105: q <= 32'b00111110010011111000010011101111 ;
        106: q <= 32'b00111110101001001011000110000000 ;
        107: q <= 32'b10111110001001100101000000110101 ;
        108: q <= 32'b00111110000111000000100001011010 ;
        109: q <= 32'b00111100010101111110001111101101 ;
        110: q <= 32'b00111101101100101100111010110101 ;
        111: q <= 32'b00111101000010000010111100010001 ;
        112: q <= 32'b10111110110011010110011101101111 ;
        113: q <= 32'b00111101101011001001111110000110 ;
        114: q <= 32'b10111110100100100111111000111111 ;
        115: q <= 32'b00111100000100111010000100111111 ;
        116: q <= 32'b00111100101111111100111010111101 ;
        117: q <= 32'b00111100000001010111011111110100 ;
        118: q <= 32'b00111110100100100111010101000000 ;
        119: q <= 32'b00111110000100111100100010010001 ;
        120: q <= 32'b10111101100100100101010100000101 ;
        121: q <= 32'b10111110011111001001100000110110 ;
        122: q <= 32'b10111110100100101010100000100001 ;
        123: q <= 32'b10111110101010100001000100000100 ;
        124: q <= 32'b00000000000000000000000000000000 ;
        125: q <= 32'b00000000000000000000000000000000 ;
        126: q <= 32'b00000000000000000000000000000000 ;
        127: q <= 32'b00000000000000000000000000000000 ;
        128: q <= 32'b00111101110000100110110111100000 ;
        129: q <= 32'b10111111000100011100111001000001 ;
        130: q <= 32'b10111110010001111010110111001011 ;
        131: q <= 32'b00111110001000110110000101110010 ;
        132: q <= 32'b00111110000100010101000000001110 ;
        133: q <= 32'b10111110101111100100101010110011 ;
        134: q <= 32'b10111101101001100010100111110100 ;
        135: q <= 32'b10111110000000111011011000101110 ;
        136: q <= 32'b00111101001100100000101000011111 ;
        137: q <= 32'b00111110011110001100010010101010 ;
        138: q <= 32'b00111101001000000101101101010111 ;
        139: q <= 32'b10111101110100010000111010011001 ;
        140: q <= 32'b00111111011010111011110011010011 ;
        141: q <= 32'b10111101110100000010100110011100 ;
        142: q <= 32'b10111111001000010101111000111001 ;
        143: q <= 32'b00111101110000110000010001010000 ;
        144: q <= 32'b10111101111011001101111010110011 ;
        145: q <= 32'b10111110001010001000110111010000 ;
        146: q <= 32'b00111111000010101101100111110010 ;
        147: q <= 32'b00111101011101011110110011100000 ;
        148: q <= 32'b10111111000000110000011001101100 ;
        149: q <= 32'b10111101011010000000100101000010 ;
        150: q <= 32'b00111111001010011000000001101110 ;
        151: q <= 32'b00111110100111001110010110010010 ;
        152: q <= 32'b10111110001000111001011110111100 ;
        153: q <= 32'b10111110000110110010101001010100 ;
        154: q <= 32'b00111110100001001100100101100000 ;
        155: q <= 32'b00111110100111001101111010111110 ;
        156: q <= 32'b00111110001011111100101001011010 ;
        157: q <= 32'b10111110101001100001110000001011 ;
        158: q <= 32'b10111110000110111011111111010111 ;
        159: q <= 32'b00111110100010111001000111100011 ;
        160: q <= 32'b00111101001101000000111110000100 ;
        161: q <= 32'b10111110010111100110011011001011 ;
        162: q <= 32'b10111110000110110101101100101010 ;
        163: q <= 32'b10111101111001101010111000001100 ;
        164: q <= 32'b00111110011010100101011111100000 ;
        165: q <= 32'b00111111010001110111000110101111 ;
        166: q <= 32'b10111110011111101100111100010000 ;
        167: q <= 32'b10111110010000000101101110110111 ;
        168: q <= 32'b10111110101000110001110000010100 ;
        169: q <= 32'b00111100100010010011100110101111 ;
        170: q <= 32'b00111110101001111110101110010101 ;
        171: q <= 32'b00111100100001001100001000111000 ;
        172: q <= 32'b00111110001000101101101000001010 ;
        173: q <= 32'b10111101111000000110110010100110 ;
        174: q <= 32'b10111110100000100001000110111110 ;
        175: q <= 32'b10111111000111100111101111000101 ;
        176: q <= 32'b10111100010100011100110000111001 ;
        177: q <= 32'b10111111001101010010010101011111 ;
        178: q <= 32'b10111110010111111010000111101001 ;
        179: q <= 32'b00111100111110110100110101000111 ;
        180: q <= 32'b10111110001111000010001111110111 ;
        181: q <= 32'b10111101001000000101110101110111 ;
        182: q <= 32'b00111110000110111110111010110010 ;
        183: q <= 32'b00111101110100011101011001001100 ;
        184: q <= 32'b10111101100100000111101010010011 ;
        185: q <= 32'b10111110100010111110101101010011 ;
        186: q <= 32'b00111110010001101100001100000011 ;
        187: q <= 32'b10111110000111000110111111100100 ;
        188: q <= 32'b00000000000000000000000000000000 ;
        189: q <= 32'b00000000000000000000000000000000 ;
        190: q <= 32'b00000000000000000000000000000000 ;
        191: q <= 32'b00000000000000000000000000000000 ;
        192: q <= 32'b00111101110101000100110100001001 ;
        193: q <= 32'b10111110101110101110101110111000 ;
        194: q <= 32'b00111111000010001001111111110011 ;
        195: q <= 32'b00111100100010101001001001001100 ;
        196: q <= 32'b00111110000001110111101111011101 ;
        197: q <= 32'b00111110101000110110000000010011 ;
        198: q <= 32'b10111101100000001101010010010110 ;
        199: q <= 32'b10111110010100111101111111110110 ;
        200: q <= 32'b00111100111001101000000010001000 ;
        201: q <= 32'b00111110001110111001110011110010 ;
        202: q <= 32'b10111111001100111110000001001011 ;
        203: q <= 32'b00111101000001111100110000011110 ;
        204: q <= 32'b00111110001110010101111001010010 ;
        205: q <= 32'b10111101100110010111111000000010 ;
        206: q <= 32'b00111101110111010101001001000111 ;
        207: q <= 32'b00111111000100100111011110110110 ;
        208: q <= 32'b00111011010010001010000110000001 ;
        209: q <= 32'b10111110001010110110111001001110 ;
        210: q <= 32'b00111101110001100101100011100110 ;
        211: q <= 32'b00111101100010000000111010000010 ;
        212: q <= 32'b00111110010110111100111001100010 ;
        213: q <= 32'b10111110000010001011101001111001 ;
        214: q <= 32'b10111101110010101101010001001101 ;
        215: q <= 32'b00111110011000100000110100010111 ;
        216: q <= 32'b10111101001101111111001110000110 ;
        217: q <= 32'b10111111001011111101100001101001 ;
        218: q <= 32'b10111110110111110100000001000010 ;
        219: q <= 32'b00111110000101011011001010110110 ;
        220: q <= 32'b00111110011001110011000010111110 ;
        221: q <= 32'b10111101110111100000011001010101 ;
        222: q <= 32'b00111101100110001110001010100110 ;
        223: q <= 32'b10111111000011110000001100010010 ;
        224: q <= 32'b10111110001001001001111111111010 ;
        225: q <= 32'b10111110100011000101001001110010 ;
        226: q <= 32'b10111110100000100011000110000101 ;
        227: q <= 32'b10111110110100101110001011101111 ;
        228: q <= 32'b00111110100000011011000011011001 ;
        229: q <= 32'b00111101000011011000101101011110 ;
        230: q <= 32'b10111110010011110100001101011010 ;
        231: q <= 32'b10111110011100101100100111111101 ;
        232: q <= 32'b10111110011111100010010110101000 ;
        233: q <= 32'b00111110000100000111000100011011 ;
        234: q <= 32'b00111110100111111111110100100101 ;
        235: q <= 32'b10111101010100110110110000000110 ;
        236: q <= 32'b00111101011110011111000100100010 ;
        237: q <= 32'b10111101101010001000011010111010 ;
        238: q <= 32'b00111110001111010111111000101101 ;
        239: q <= 32'b10111111000011100111000100110001 ;
        240: q <= 32'b00111110011110100100101100100010 ;
        241: q <= 32'b00111101110010101000000000110110 ;
        242: q <= 32'b10111110001110010101110010011011 ;
        243: q <= 32'b00111111010110001101100101000100 ;
        244: q <= 32'b10111100110010111111000111011110 ;
        245: q <= 32'b00111111000001011000100100101001 ;
        246: q <= 32'b00111110011010101011011110100110 ;
        247: q <= 32'b00111110001010001011001111000001 ;
        248: q <= 32'b00111110000101100101101001100111 ;
        249: q <= 32'b10111110100001011101110110110101 ;
        250: q <= 32'b00111110110111110001001011101000 ;
        251: q <= 32'b10111110010001100010110101000010 ;
        252: q <= 32'b00000000000000000000000000000000 ;
        253: q <= 32'b00000000000000000000000000000000 ;
        254: q <= 32'b00000000000000000000000000000000 ;
        255: q <= 32'b00000000000000000000000000000000 ;
        256: q <= 32'b00000000000000000000000000000000 ;
        257: q <= 32'b00000000000000000000000000000000 ;
        258: q <= 32'b00000000000000000000000000000000 ;
        259: q <= 32'b00000000000000000000000000000000 ;
        260: q <= 32'b00000000000000000000000000000000 ;
        261: q <= 32'b00000000000000000000000000000000 ;
        262: q <= 32'b00000000000000000000000000000000 ;
        263: q <= 32'b00000000000000000000000000000000 ;
        264: q <= 32'b00000000000000000000000000000000 ;
        265: q <= 32'b00000000000000000000000000000000 ;
        266: q <= 32'b00000000000000000000000000000000 ;
        267: q <= 32'b00000000000000000000000000000000 ;
        268: q <= 32'b00000000000000000000000000000000 ;
        269: q <= 32'b00000000000000000000000000000000 ;
        270: q <= 32'b00000000000000000000000000000000 ;
        271: q <= 32'b00000000000000000000000000000000 ;
        272: q <= 32'b00000000000000000000000000000000 ;
        273: q <= 32'b00000000000000000000000000000000 ;
        274: q <= 32'b00000000000000000000000000000000 ;
        275: q <= 32'b00000000000000000000000000000000 ;
        276: q <= 32'b00000000000000000000000000000000 ;
        277: q <= 32'b00000000000000000000000000000000 ;
        278: q <= 32'b00000000000000000000000000000000 ;
        279: q <= 32'b00000000000000000000000000000000 ;
        280: q <= 32'b00000000000000000000000000000000 ;
        281: q <= 32'b00000000000000000000000000000000 ;
        282: q <= 32'b00000000000000000000000000000000 ;
        283: q <= 32'b00000000000000000000000000000000 ;
        284: q <= 32'b00000000000000000000000000000000 ;
        285: q <= 32'b00000000000000000000000000000000 ;
        286: q <= 32'b00000000000000000000000000000000 ;
        287: q <= 32'b00000000000000000000000000000000 ;
        288: q <= 32'b00000000000000000000000000000000 ;
        289: q <= 32'b00000000000000000000000000000000 ;
        290: q <= 32'b00000000000000000000000000000000 ;
        291: q <= 32'b00000000000000000000000000000000 ;
        292: q <= 32'b00000000000000000000000000000000 ;
        293: q <= 32'b00000000000000000000000000000000 ;
        294: q <= 32'b00000000000000000000000000000000 ;
        295: q <= 32'b00000000000000000000000000000000 ;
        296: q <= 32'b00000000000000000000000000000000 ;
        297: q <= 32'b00000000000000000000000000000000 ;
        298: q <= 32'b00000000000000000000000000000000 ;
        299: q <= 32'b00000000000000000000000000000000 ;
        300: q <= 32'b00000000000000000000000000000000 ;
        301: q <= 32'b00000000000000000000000000000000 ;
        302: q <= 32'b00000000000000000000000000000000 ;
        303: q <= 32'b00000000000000000000000000000000 ;
        304: q <= 32'b00000000000000000000000000000000 ;
        305: q <= 32'b00000000000000000000000000000000 ;
        306: q <= 32'b00000000000000000000000000000000 ;
        307: q <= 32'b00000000000000000000000000000000 ;
        308: q <= 32'b00000000000000000000000000000000 ;
        309: q <= 32'b00000000000000000000000000000000 ;
        310: q <= 32'b00000000000000000000000000000000 ;
        311: q <= 32'b00000000000000000000000000000000 ;
        312: q <= 32'b00000000000000000000000000000000 ;
        313: q <= 32'b00000000000000000000000000000000 ;
        314: q <= 32'b00000000000000000000000000000000 ;
        315: q <= 32'b00000000000000000000000000000000 ;
        316: q <= 32'b00000000000000000000000000000000 ;
        317: q <= 32'b00000000000000000000000000000000 ;
        318: q <= 32'b00000000000000000000000000000000 ;
        319: q <= 32'b00000000000000000000000000000000 ;
        320: q <= 32'b00000000000000000000000000000000 ;
        321: q <= 32'b00000000000000000000000000000000 ;
        322: q <= 32'b00000000000000000000000000000000 ;
        323: q <= 32'b00000000000000000000000000000000 ;
        324: q <= 32'b00000000000000000000000000000000 ;
        325: q <= 32'b00000000000000000000000000000000 ;
        326: q <= 32'b00000000000000000000000000000000 ;
        327: q <= 32'b00000000000000000000000000000000 ;
        328: q <= 32'b00000000000000000000000000000000 ;
        329: q <= 32'b00000000000000000000000000000000 ;
        330: q <= 32'b00000000000000000000000000000000 ;
        331: q <= 32'b00000000000000000000000000000000 ;
        332: q <= 32'b00000000000000000000000000000000 ;
        333: q <= 32'b00000000000000000000000000000000 ;
        334: q <= 32'b00000000000000000000000000000000 ;
        335: q <= 32'b00000000000000000000000000000000 ;
        336: q <= 32'b00000000000000000000000000000000 ;
        337: q <= 32'b00000000000000000000000000000000 ;
        338: q <= 32'b00000000000000000000000000000000 ;
        339: q <= 32'b00000000000000000000000000000000 ;
        340: q <= 32'b00000000000000000000000000000000 ;
        341: q <= 32'b00000000000000000000000000000000 ;
        342: q <= 32'b00000000000000000000000000000000 ;
        343: q <= 32'b00000000000000000000000000000000 ;
        344: q <= 32'b00000000000000000000000000000000 ;
        345: q <= 32'b00000000000000000000000000000000 ;
        346: q <= 32'b00000000000000000000000000000000 ;
        347: q <= 32'b00000000000000000000000000000000 ;
        348: q <= 32'b00000000000000000000000000000000 ;
        349: q <= 32'b00000000000000000000000000000000 ;
        350: q <= 32'b00000000000000000000000000000000 ;
        351: q <= 32'b00000000000000000000000000000000 ;
        352: q <= 32'b00000000000000000000000000000000 ;
        353: q <= 32'b00000000000000000000000000000000 ;
        354: q <= 32'b00000000000000000000000000000000 ;
        355: q <= 32'b00000000000000000000000000000000 ;
        356: q <= 32'b00000000000000000000000000000000 ;
        357: q <= 32'b00000000000000000000000000000000 ;
        358: q <= 32'b00000000000000000000000000000000 ;
        359: q <= 32'b00000000000000000000000000000000 ;
        360: q <= 32'b00000000000000000000000000000000 ;
        361: q <= 32'b00000000000000000000000000000000 ;
        362: q <= 32'b00000000000000000000000000000000 ;
        363: q <= 32'b00000000000000000000000000000000 ;
        364: q <= 32'b00000000000000000000000000000000 ;
        365: q <= 32'b00000000000000000000000000000000 ;
        366: q <= 32'b00000000000000000000000000000000 ;
        367: q <= 32'b00000000000000000000000000000000 ;
        368: q <= 32'b00000000000000000000000000000000 ;
        369: q <= 32'b00000000000000000000000000000000 ;
        370: q <= 32'b00000000000000000000000000000000 ;
        371: q <= 32'b00000000000000000000000000000000 ;
        372: q <= 32'b00000000000000000000000000000000 ;
        373: q <= 32'b00000000000000000000000000000000 ;
        374: q <= 32'b00000000000000000000000000000000 ;
        375: q <= 32'b00000000000000000000000000000000 ;
        376: q <= 32'b00000000000000000000000000000000 ;
        377: q <= 32'b00000000000000000000000000000000 ;
        378: q <= 32'b00000000000000000000000000000000 ;
        379: q <= 32'b00000000000000000000000000000000 ;
        380: q <= 32'b00000000000000000000000000000000 ;
        381: q <= 32'b00000000000000000000000000000000 ;
        382: q <= 32'b00000000000000000000000000000000 ;
        383: q <= 32'b00000000000000000000000000000000 ;
        384: q <= 32'b00000000000000000000000000000000 ;
        385: q <= 32'b00000000000000000000000000000000 ;
        386: q <= 32'b00000000000000000000000000000000 ;
        387: q <= 32'b00000000000000000000000000000000 ;
        388: q <= 32'b00000000000000000000000000000000 ;
        389: q <= 32'b00000000000000000000000000000000 ;
        390: q <= 32'b00000000000000000000000000000000 ;
        391: q <= 32'b00000000000000000000000000000000 ;
        392: q <= 32'b00000000000000000000000000000000 ;
        393: q <= 32'b00000000000000000000000000000000 ;
        394: q <= 32'b00000000000000000000000000000000 ;
        395: q <= 32'b00000000000000000000000000000000 ;
        396: q <= 32'b00000000000000000000000000000000 ;
        397: q <= 32'b00000000000000000000000000000000 ;
        398: q <= 32'b00000000000000000000000000000000 ;
        399: q <= 32'b00000000000000000000000000000000 ;
        400: q <= 32'b00000000000000000000000000000000 ;
        401: q <= 32'b00000000000000000000000000000000 ;
        402: q <= 32'b00000000000000000000000000000000 ;
        403: q <= 32'b00000000000000000000000000000000 ;
        404: q <= 32'b00000000000000000000000000000000 ;
        405: q <= 32'b00000000000000000000000000000000 ;
        406: q <= 32'b00000000000000000000000000000000 ;
        407: q <= 32'b00000000000000000000000000000000 ;
        408: q <= 32'b00000000000000000000000000000000 ;
        409: q <= 32'b00000000000000000000000000000000 ;
        410: q <= 32'b00000000000000000000000000000000 ;
        411: q <= 32'b00000000000000000000000000000000 ;
        412: q <= 32'b00000000000000000000000000000000 ;
        413: q <= 32'b00000000000000000000000000000000 ;
        414: q <= 32'b00000000000000000000000000000000 ;
        415: q <= 32'b00000000000000000000000000000000 ;
        416: q <= 32'b00000000000000000000000000000000 ;
        417: q <= 32'b00000000000000000000000000000000 ;
        418: q <= 32'b00000000000000000000000000000000 ;
        419: q <= 32'b00000000000000000000000000000000 ;
        420: q <= 32'b00000000000000000000000000000000 ;
        421: q <= 32'b00000000000000000000000000000000 ;
        422: q <= 32'b00000000000000000000000000000000 ;
        423: q <= 32'b00000000000000000000000000000000 ;
        424: q <= 32'b00000000000000000000000000000000 ;
        425: q <= 32'b00000000000000000000000000000000 ;
        426: q <= 32'b00000000000000000000000000000000 ;
        427: q <= 32'b00000000000000000000000000000000 ;
        428: q <= 32'b00000000000000000000000000000000 ;
        429: q <= 32'b00000000000000000000000000000000 ;
        430: q <= 32'b00000000000000000000000000000000 ;
        431: q <= 32'b00000000000000000000000000000000 ;
        432: q <= 32'b00000000000000000000000000000000 ;
        433: q <= 32'b00000000000000000000000000000000 ;
        434: q <= 32'b00000000000000000000000000000000 ;
        435: q <= 32'b00000000000000000000000000000000 ;
        436: q <= 32'b00000000000000000000000000000000 ;
        437: q <= 32'b00000000000000000000000000000000 ;
        438: q <= 32'b00000000000000000000000000000000 ;
        439: q <= 32'b00000000000000000000000000000000 ;
        440: q <= 32'b00000000000000000000000000000000 ;
        441: q <= 32'b00000000000000000000000000000000 ;
        442: q <= 32'b00000000000000000000000000000000 ;
        443: q <= 32'b00000000000000000000000000000000 ;
        444: q <= 32'b00000000000000000000000000000000 ;
        445: q <= 32'b00000000000000000000000000000000 ;
        446: q <= 32'b00000000000000000000000000000000 ;
        447: q <= 32'b00000000000000000000000000000000 ;
        448: q <= 32'b00000000000000000000000000000000 ;
        449: q <= 32'b00000000000000000000000000000000 ;
        450: q <= 32'b00000000000000000000000000000000 ;
        451: q <= 32'b00000000000000000000000000000000 ;
        452: q <= 32'b00000000000000000000000000000000 ;
        453: q <= 32'b00000000000000000000000000000000 ;
        454: q <= 32'b00000000000000000000000000000000 ;
        455: q <= 32'b00000000000000000000000000000000 ;
        456: q <= 32'b00000000000000000000000000000000 ;
        457: q <= 32'b00000000000000000000000000000000 ;
        458: q <= 32'b00000000000000000000000000000000 ;
        459: q <= 32'b00000000000000000000000000000000 ;
        460: q <= 32'b00000000000000000000000000000000 ;
        461: q <= 32'b00000000000000000000000000000000 ;
        462: q <= 32'b00000000000000000000000000000000 ;
        463: q <= 32'b00000000000000000000000000000000 ;
        464: q <= 32'b00000000000000000000000000000000 ;
        465: q <= 32'b00000000000000000000000000000000 ;
        466: q <= 32'b00000000000000000000000000000000 ;
        467: q <= 32'b00000000000000000000000000000000 ;
        468: q <= 32'b00000000000000000000000000000000 ;
        469: q <= 32'b00000000000000000000000000000000 ;
        470: q <= 32'b00000000000000000000000000000000 ;
        471: q <= 32'b00000000000000000000000000000000 ;
        472: q <= 32'b00000000000000000000000000000000 ;
        473: q <= 32'b00000000000000000000000000000000 ;
        474: q <= 32'b00000000000000000000000000000000 ;
        475: q <= 32'b00000000000000000000000000000000 ;
        476: q <= 32'b00000000000000000000000000000000 ;
        477: q <= 32'b00000000000000000000000000000000 ;
        478: q <= 32'b00000000000000000000000000000000 ;
        479: q <= 32'b00000000000000000000000000000000 ;
        480: q <= 32'b00000000000000000000000000000000 ;
        481: q <= 32'b00000000000000000000000000000000 ;
        482: q <= 32'b00000000000000000000000000000000 ;
        483: q <= 32'b00000000000000000000000000000000 ;
        484: q <= 32'b00000000000000000000000000000000 ;
        485: q <= 32'b00000000000000000000000000000000 ;
        486: q <= 32'b00000000000000000000000000000000 ;
        487: q <= 32'b00000000000000000000000000000000 ;
        488: q <= 32'b00000000000000000000000000000000 ;
        489: q <= 32'b00000000000000000000000000000000 ;
        490: q <= 32'b00000000000000000000000000000000 ;
        491: q <= 32'b00000000000000000000000000000000 ;
        492: q <= 32'b00000000000000000000000000000000 ;
        493: q <= 32'b00000000000000000000000000000000 ;
        494: q <= 32'b00000000000000000000000000000000 ;
        495: q <= 32'b00000000000000000000000000000000 ;
        496: q <= 32'b00000000000000000000000000000000 ;
        497: q <= 32'b00000000000000000000000000000000 ;
        498: q <= 32'b00000000000000000000000000000000 ;
        499: q <= 32'b00000000000000000000000000000000 ;
        500: q <= 32'b00000000000000000000000000000000 ;
        501: q <= 32'b00000000000000000000000000000000 ;
        502: q <= 32'b00000000000000000000000000000000 ;
        503: q <= 32'b00000000000000000000000000000000 ;
        504: q <= 32'b00000000000000000000000000000000 ;
        505: q <= 32'b00000000000000000000000000000000 ;
        506: q <= 32'b00000000000000000000000000000000 ;
        507: q <= 32'b00000000000000000000000000000000 ;
        508: q <= 32'b00000000000000000000000000000000 ;
        509: q <= 32'b00000000000000000000000000000000 ;
        510: q <= 32'b00000000000000000000000000000000 ;
        511: q <= 32'b00000000000000000000000000000000 ;
        512: q <= 32'b00000000000000000000000000000000 ;
        513: q <= 32'b00000000000000000000000000000000 ;
        514: q <= 32'b00000000000000000000000000000000 ;
        515: q <= 32'b00000000000000000000000000000000 ;
        516: q <= 32'b00000000000000000000000000000000 ;
        517: q <= 32'b00000000000000000000000000000000 ;
        518: q <= 32'b00000000000000000000000000000000 ;
        519: q <= 32'b00000000000000000000000000000000 ;
        520: q <= 32'b00000000000000000000000000000000 ;
        521: q <= 32'b00000000000000000000000000000000 ;
        522: q <= 32'b00000000000000000000000000000000 ;
        523: q <= 32'b00000000000000000000000000000000 ;
        524: q <= 32'b00000000000000000000000000000000 ;
        525: q <= 32'b00000000000000000000000000000000 ;
        526: q <= 32'b00000000000000000000000000000000 ;
        527: q <= 32'b00000000000000000000000000000000 ;
        528: q <= 32'b00000000000000000000000000000000 ;
        529: q <= 32'b00000000000000000000000000000000 ;
        530: q <= 32'b00000000000000000000000000000000 ;
        531: q <= 32'b00000000000000000000000000000000 ;
        532: q <= 32'b00000000000000000000000000000000 ;
        533: q <= 32'b00000000000000000000000000000000 ;
        534: q <= 32'b00000000000000000000000000000000 ;
        535: q <= 32'b00000000000000000000000000000000 ;
        536: q <= 32'b00000000000000000000000000000000 ;
        537: q <= 32'b00000000000000000000000000000000 ;
        538: q <= 32'b00000000000000000000000000000000 ;
        539: q <= 32'b00000000000000000000000000000000 ;
        540: q <= 32'b00000000000000000000000000000000 ;
        541: q <= 32'b00000000000000000000000000000000 ;
        542: q <= 32'b00000000000000000000000000000000 ;
        543: q <= 32'b00000000000000000000000000000000 ;
        544: q <= 32'b00000000000000000000000000000000 ;
        545: q <= 32'b00000000000000000000000000000000 ;
        546: q <= 32'b00000000000000000000000000000000 ;
        547: q <= 32'b00000000000000000000000000000000 ;
        548: q <= 32'b00000000000000000000000000000000 ;
        549: q <= 32'b00000000000000000000000000000000 ;
        550: q <= 32'b00000000000000000000000000000000 ;
        551: q <= 32'b00000000000000000000000000000000 ;
        552: q <= 32'b00000000000000000000000000000000 ;
        553: q <= 32'b00000000000000000000000000000000 ;
        554: q <= 32'b00000000000000000000000000000000 ;
        555: q <= 32'b00000000000000000000000000000000 ;
        556: q <= 32'b00000000000000000000000000000000 ;
        557: q <= 32'b00000000000000000000000000000000 ;
        558: q <= 32'b00000000000000000000000000000000 ;
        559: q <= 32'b00000000000000000000000000000000 ;
        560: q <= 32'b00000000000000000000000000000000 ;
        561: q <= 32'b00000000000000000000000000000000 ;
        562: q <= 32'b00000000000000000000000000000000 ;
        563: q <= 32'b00000000000000000000000000000000 ;
        564: q <= 32'b00000000000000000000000000000000 ;
        565: q <= 32'b00000000000000000000000000000000 ;
        566: q <= 32'b00000000000000000000000000000000 ;
        567: q <= 32'b00000000000000000000000000000000 ;
        568: q <= 32'b00000000000000000000000000000000 ;
        569: q <= 32'b00000000000000000000000000000000 ;
        570: q <= 32'b00000000000000000000000000000000 ;
        571: q <= 32'b00000000000000000000000000000000 ;
        572: q <= 32'b00000000000000000000000000000000 ;
        573: q <= 32'b00000000000000000000000000000000 ;
        574: q <= 32'b00000000000000000000000000000000 ;
        575: q <= 32'b00000000000000000000000000000000 ;
        576: q <= 32'b00000000000000000000000000000000 ;
        577: q <= 32'b00000000000000000000000000000000 ;
        578: q <= 32'b00000000000000000000000000000000 ;
        579: q <= 32'b00000000000000000000000000000000 ;
        580: q <= 32'b00000000000000000000000000000000 ;
        581: q <= 32'b00000000000000000000000000000000 ;
        582: q <= 32'b00000000000000000000000000000000 ;
        583: q <= 32'b00000000000000000000000000000000 ;
        584: q <= 32'b00000000000000000000000000000000 ;
        585: q <= 32'b00000000000000000000000000000000 ;
        586: q <= 32'b00000000000000000000000000000000 ;
        587: q <= 32'b00000000000000000000000000000000 ;
        588: q <= 32'b00000000000000000000000000000000 ;
        589: q <= 32'b00000000000000000000000000000000 ;
        590: q <= 32'b00000000000000000000000000000000 ;
        591: q <= 32'b00000000000000000000000000000000 ;
        592: q <= 32'b00000000000000000000000000000000 ;
        593: q <= 32'b00000000000000000000000000000000 ;
        594: q <= 32'b00000000000000000000000000000000 ;
        595: q <= 32'b00000000000000000000000000000000 ;
        596: q <= 32'b00000000000000000000000000000000 ;
        597: q <= 32'b00000000000000000000000000000000 ;
        598: q <= 32'b00000000000000000000000000000000 ;
        599: q <= 32'b00000000000000000000000000000000 ;
        600: q <= 32'b00000000000000000000000000000000 ;
        601: q <= 32'b00000000000000000000000000000000 ;
        602: q <= 32'b00000000000000000000000000000000 ;
        603: q <= 32'b00000000000000000000000000000000 ;
        604: q <= 32'b00000000000000000000000000000000 ;
        605: q <= 32'b00000000000000000000000000000000 ;
        606: q <= 32'b00000000000000000000000000000000 ;
        607: q <= 32'b00000000000000000000000000000000 ;
        608: q <= 32'b00000000000000000000000000000000 ;
        609: q <= 32'b00000000000000000000000000000000 ;
        610: q <= 32'b00000000000000000000000000000000 ;
        611: q <= 32'b00000000000000000000000000000000 ;
        612: q <= 32'b00000000000000000000000000000000 ;
        613: q <= 32'b00000000000000000000000000000000 ;
        614: q <= 32'b00000000000000000000000000000000 ;
        615: q <= 32'b00000000000000000000000000000000 ;
        616: q <= 32'b00000000000000000000000000000000 ;
        617: q <= 32'b00000000000000000000000000000000 ;
        618: q <= 32'b00000000000000000000000000000000 ;
        619: q <= 32'b00000000000000000000000000000000 ;
        620: q <= 32'b00000000000000000000000000000000 ;
        621: q <= 32'b00000000000000000000000000000000 ;
        622: q <= 32'b00000000000000000000000000000000 ;
        623: q <= 32'b00000000000000000000000000000000 ;
        624: q <= 32'b00000000000000000000000000000000 ;
        625: q <= 32'b00000000000000000000000000000000 ;
        626: q <= 32'b00000000000000000000000000000000 ;
        627: q <= 32'b00000000000000000000000000000000 ;
        628: q <= 32'b00000000000000000000000000000000 ;
        629: q <= 32'b00000000000000000000000000000000 ;
        630: q <= 32'b00000000000000000000000000000000 ;
        631: q <= 32'b00000000000000000000000000000000 ;
        632: q <= 32'b00000000000000000000000000000000 ;
        633: q <= 32'b00000000000000000000000000000000 ;
        634: q <= 32'b00000000000000000000000000000000 ;
        635: q <= 32'b00000000000000000000000000000000 ;
        636: q <= 32'b00000000000000000000000000000000 ;
        637: q <= 32'b00000000000000000000000000000000 ;
        638: q <= 32'b00000000000000000000000000000000 ;
        639: q <= 32'b00000000000000000000000000000000 ;
        640: q <= 32'b00000000000000000000000000000000 ;
        641: q <= 32'b00000000000000000000000000000000 ;
        642: q <= 32'b00000000000000000000000000000000 ;
        643: q <= 32'b00000000000000000000000000000000 ;
        644: q <= 32'b00000000000000000000000000000000 ;
        645: q <= 32'b00000000000000000000000000000000 ;
        646: q <= 32'b00000000000000000000000000000000 ;
        647: q <= 32'b00000000000000000000000000000000 ;
        648: q <= 32'b00000000000000000000000000000000 ;
        649: q <= 32'b00000000000000000000000000000000 ;
        650: q <= 32'b00000000000000000000000000000000 ;
        651: q <= 32'b00000000000000000000000000000000 ;
        652: q <= 32'b00000000000000000000000000000000 ;
        653: q <= 32'b00000000000000000000000000000000 ;
        654: q <= 32'b00000000000000000000000000000000 ;
        655: q <= 32'b00000000000000000000000000000000 ;
        656: q <= 32'b00000000000000000000000000000000 ;
        657: q <= 32'b00000000000000000000000000000000 ;
        658: q <= 32'b00000000000000000000000000000000 ;
        659: q <= 32'b00000000000000000000000000000000 ;
        660: q <= 32'b00000000000000000000000000000000 ;
        661: q <= 32'b00000000000000000000000000000000 ;
        662: q <= 32'b00000000000000000000000000000000 ;
        663: q <= 32'b00000000000000000000000000000000 ;
        664: q <= 32'b00000000000000000000000000000000 ;
        665: q <= 32'b00000000000000000000000000000000 ;
        666: q <= 32'b00000000000000000000000000000000 ;
        667: q <= 32'b00000000000000000000000000000000 ;
        668: q <= 32'b00000000000000000000000000000000 ;
        669: q <= 32'b00000000000000000000000000000000 ;
        670: q <= 32'b00000000000000000000000000000000 ;
        671: q <= 32'b00000000000000000000000000000000 ;
        672: q <= 32'b00000000000000000000000000000000 ;
        673: q <= 32'b00000000000000000000000000000000 ;
        674: q <= 32'b00000000000000000000000000000000 ;
        675: q <= 32'b00000000000000000000000000000000 ;
        676: q <= 32'b00000000000000000000000000000000 ;
        677: q <= 32'b00000000000000000000000000000000 ;
        678: q <= 32'b00000000000000000000000000000000 ;
        679: q <= 32'b00000000000000000000000000000000 ;
        680: q <= 32'b00000000000000000000000000000000 ;
        681: q <= 32'b00000000000000000000000000000000 ;
        682: q <= 32'b00000000000000000000000000000000 ;
        683: q <= 32'b00000000000000000000000000000000 ;
        684: q <= 32'b00000000000000000000000000000000 ;
        685: q <= 32'b00000000000000000000000000000000 ;
        686: q <= 32'b00000000000000000000000000000000 ;
        687: q <= 32'b00000000000000000000000000000000 ;
        688: q <= 32'b00000000000000000000000000000000 ;
        689: q <= 32'b00000000000000000000000000000000 ;
        690: q <= 32'b00000000000000000000000000000000 ;
        691: q <= 32'b00000000000000000000000000000000 ;
        692: q <= 32'b00000000000000000000000000000000 ;
        693: q <= 32'b00000000000000000000000000000000 ;
        694: q <= 32'b00000000000000000000000000000000 ;
        695: q <= 32'b00000000000000000000000000000000 ;
        696: q <= 32'b00000000000000000000000000000000 ;
        697: q <= 32'b00000000000000000000000000000000 ;
        698: q <= 32'b00000000000000000000000000000000 ;
        699: q <= 32'b00000000000000000000000000000000 ;
        700: q <= 32'b00000000000000000000000000000000 ;
        701: q <= 32'b00000000000000000000000000000000 ;
        702: q <= 32'b00000000000000000000000000000000 ;
        703: q <= 32'b00000000000000000000000000000000 ;
        704: q <= 32'b00000000000000000000000000000000 ;
        705: q <= 32'b00000000000000000000000000000000 ;
        706: q <= 32'b00000000000000000000000000000000 ;
        707: q <= 32'b00000000000000000000000000000000 ;
        708: q <= 32'b00000000000000000000000000000000 ;
        709: q <= 32'b00000000000000000000000000000000 ;
        710: q <= 32'b00000000000000000000000000000000 ;
        711: q <= 32'b00000000000000000000000000000000 ;
        712: q <= 32'b00000000000000000000000000000000 ;
        713: q <= 32'b00000000000000000000000000000000 ;
        714: q <= 32'b00000000000000000000000000000000 ;
        715: q <= 32'b00000000000000000000000000000000 ;
        716: q <= 32'b00000000000000000000000000000000 ;
        717: q <= 32'b00000000000000000000000000000000 ;
        718: q <= 32'b00000000000000000000000000000000 ;
        719: q <= 32'b00000000000000000000000000000000 ;
        720: q <= 32'b00000000000000000000000000000000 ;
        721: q <= 32'b00000000000000000000000000000000 ;
        722: q <= 32'b00000000000000000000000000000000 ;
        723: q <= 32'b00000000000000000000000000000000 ;
        724: q <= 32'b00000000000000000000000000000000 ;
        725: q <= 32'b00000000000000000000000000000000 ;
        726: q <= 32'b00000000000000000000000000000000 ;
        727: q <= 32'b00000000000000000000000000000000 ;
        728: q <= 32'b00000000000000000000000000000000 ;
        729: q <= 32'b00000000000000000000000000000000 ;
        730: q <= 32'b00000000000000000000000000000000 ;
        731: q <= 32'b00000000000000000000000000000000 ;
        732: q <= 32'b00000000000000000000000000000000 ;
        733: q <= 32'b00000000000000000000000000000000 ;
        734: q <= 32'b00000000000000000000000000000000 ;
        735: q <= 32'b00000000000000000000000000000000 ;
        736: q <= 32'b00000000000000000000000000000000 ;
        737: q <= 32'b00000000000000000000000000000000 ;
        738: q <= 32'b00000000000000000000000000000000 ;
        739: q <= 32'b00000000000000000000000000000000 ;
        740: q <= 32'b00000000000000000000000000000000 ;
        741: q <= 32'b00000000000000000000000000000000 ;
        742: q <= 32'b00000000000000000000000000000000 ;
        743: q <= 32'b00000000000000000000000000000000 ;
        744: q <= 32'b00000000000000000000000000000000 ;
        745: q <= 32'b00000000000000000000000000000000 ;
        746: q <= 32'b00000000000000000000000000000000 ;
        747: q <= 32'b00000000000000000000000000000000 ;
        748: q <= 32'b00000000000000000000000000000000 ;
        749: q <= 32'b00000000000000000000000000000000 ;
        750: q <= 32'b00000000000000000000000000000000 ;
        751: q <= 32'b00000000000000000000000000000000 ;
        752: q <= 32'b00000000000000000000000000000000 ;
        753: q <= 32'b00000000000000000000000000000000 ;
        754: q <= 32'b00000000000000000000000000000000 ;
        755: q <= 32'b00000000000000000000000000000000 ;
        756: q <= 32'b00000000000000000000000000000000 ;
        757: q <= 32'b00000000000000000000000000000000 ;
        758: q <= 32'b00000000000000000000000000000000 ;
        759: q <= 32'b00000000000000000000000000000000 ;
        760: q <= 32'b00000000000000000000000000000000 ;
        761: q <= 32'b00000000000000000000000000000000 ;
        762: q <= 32'b00000000000000000000000000000000 ;
        763: q <= 32'b00000000000000000000000000000000 ;
        764: q <= 32'b00000000000000000000000000000000 ;
        765: q <= 32'b00000000000000000000000000000000 ;
        766: q <= 32'b00000000000000000000000000000000 ;
        767: q <= 32'b00000000000000000000000000000000 ;
        768: q <= 32'b00000000000000000000000000000000 ;
        769: q <= 32'b00000000000000000000000000000000 ;
        770: q <= 32'b00000000000000000000000000000000 ;
        771: q <= 32'b00000000000000000000000000000000 ;
        772: q <= 32'b00000000000000000000000000000000 ;
        773: q <= 32'b00000000000000000000000000000000 ;
        774: q <= 32'b00000000000000000000000000000000 ;
        775: q <= 32'b00000000000000000000000000000000 ;
        776: q <= 32'b00000000000000000000000000000000 ;
        777: q <= 32'b00000000000000000000000000000000 ;
        778: q <= 32'b00000000000000000000000000000000 ;
        779: q <= 32'b00000000000000000000000000000000 ;
        780: q <= 32'b00000000000000000000000000000000 ;
        781: q <= 32'b00000000000000000000000000000000 ;
        782: q <= 32'b00000000000000000000000000000000 ;
        783: q <= 32'b00000000000000000000000000000000 ;
        784: q <= 32'b00000000000000000000000000000000 ;
        785: q <= 32'b00000000000000000000000000000000 ;
        786: q <= 32'b00000000000000000000000000000000 ;
        787: q <= 32'b00000000000000000000000000000000 ;
        788: q <= 32'b00000000000000000000000000000000 ;
        789: q <= 32'b00000000000000000000000000000000 ;
        790: q <= 32'b00000000000000000000000000000000 ;
        791: q <= 32'b00000000000000000000000000000000 ;
        792: q <= 32'b00000000000000000000000000000000 ;
        793: q <= 32'b00000000000000000000000000000000 ;
        794: q <= 32'b00000000000000000000000000000000 ;
        795: q <= 32'b00000000000000000000000000000000 ;
        796: q <= 32'b00000000000000000000000000000000 ;
        797: q <= 32'b00000000000000000000000000000000 ;
        798: q <= 32'b00000000000000000000000000000000 ;
        799: q <= 32'b00000000000000000000000000000000 ;
        800: q <= 32'b00000000000000000000000000000000 ;
        801: q <= 32'b00000000000000000000000000000000 ;
        802: q <= 32'b00000000000000000000000000000000 ;
        803: q <= 32'b00000000000000000000000000000000 ;
        804: q <= 32'b00000000000000000000000000000000 ;
        805: q <= 32'b00000000000000000000000000000000 ;
        806: q <= 32'b00000000000000000000000000000000 ;
        807: q <= 32'b00000000000000000000000000000000 ;
        808: q <= 32'b00000000000000000000000000000000 ;
        809: q <= 32'b00000000000000000000000000000000 ;
        810: q <= 32'b00000000000000000000000000000000 ;
        811: q <= 32'b00000000000000000000000000000000 ;
        812: q <= 32'b00000000000000000000000000000000 ;
        813: q <= 32'b00000000000000000000000000000000 ;
        814: q <= 32'b00000000000000000000000000000000 ;
        815: q <= 32'b00000000000000000000000000000000 ;
        816: q <= 32'b00000000000000000000000000000000 ;
        817: q <= 32'b00000000000000000000000000000000 ;
        818: q <= 32'b00000000000000000000000000000000 ;
        819: q <= 32'b00000000000000000000000000000000 ;
        820: q <= 32'b00000000000000000000000000000000 ;
        821: q <= 32'b00000000000000000000000000000000 ;
        822: q <= 32'b00000000000000000000000000000000 ;
        823: q <= 32'b00000000000000000000000000000000 ;
        824: q <= 32'b00000000000000000000000000000000 ;
        825: q <= 32'b00000000000000000000000000000000 ;
        826: q <= 32'b00000000000000000000000000000000 ;
        827: q <= 32'b00000000000000000000000000000000 ;
        828: q <= 32'b00000000000000000000000000000000 ;
        829: q <= 32'b00000000000000000000000000000000 ;
        830: q <= 32'b00000000000000000000000000000000 ;
        831: q <= 32'b00000000000000000000000000000000 ;
        832: q <= 32'b00000000000000000000000000000000 ;
        833: q <= 32'b00000000000000000000000000000000 ;
        834: q <= 32'b00000000000000000000000000000000 ;
        835: q <= 32'b00000000000000000000000000000000 ;
        836: q <= 32'b00000000000000000000000000000000 ;
        837: q <= 32'b00000000000000000000000000000000 ;
        838: q <= 32'b00000000000000000000000000000000 ;
        839: q <= 32'b00000000000000000000000000000000 ;
        840: q <= 32'b00000000000000000000000000000000 ;
        841: q <= 32'b00000000000000000000000000000000 ;
        842: q <= 32'b00000000000000000000000000000000 ;
        843: q <= 32'b00000000000000000000000000000000 ;
        844: q <= 32'b00000000000000000000000000000000 ;
        845: q <= 32'b00000000000000000000000000000000 ;
        846: q <= 32'b00000000000000000000000000000000 ;
        847: q <= 32'b00000000000000000000000000000000 ;
        848: q <= 32'b00000000000000000000000000000000 ;
        849: q <= 32'b00000000000000000000000000000000 ;
        850: q <= 32'b00000000000000000000000000000000 ;
        851: q <= 32'b00000000000000000000000000000000 ;
        852: q <= 32'b00000000000000000000000000000000 ;
        853: q <= 32'b00000000000000000000000000000000 ;
        854: q <= 32'b00000000000000000000000000000000 ;
        855: q <= 32'b00000000000000000000000000000000 ;
        856: q <= 32'b00000000000000000000000000000000 ;
        857: q <= 32'b00000000000000000000000000000000 ;
        858: q <= 32'b00000000000000000000000000000000 ;
        859: q <= 32'b00000000000000000000000000000000 ;
        860: q <= 32'b00000000000000000000000000000000 ;
        861: q <= 32'b00000000000000000000000000000000 ;
        862: q <= 32'b00000000000000000000000000000000 ;
        863: q <= 32'b00000000000000000000000000000000 ;
        864: q <= 32'b00000000000000000000000000000000 ;
        865: q <= 32'b00000000000000000000000000000000 ;
        866: q <= 32'b00000000000000000000000000000000 ;
        867: q <= 32'b00000000000000000000000000000000 ;
        868: q <= 32'b00000000000000000000000000000000 ;
        869: q <= 32'b00000000000000000000000000000000 ;
        870: q <= 32'b00000000000000000000000000000000 ;
        871: q <= 32'b00000000000000000000000000000000 ;
        872: q <= 32'b00000000000000000000000000000000 ;
        873: q <= 32'b00000000000000000000000000000000 ;
        874: q <= 32'b00000000000000000000000000000000 ;
        875: q <= 32'b00000000000000000000000000000000 ;
        876: q <= 32'b00000000000000000000000000000000 ;
        877: q <= 32'b00000000000000000000000000000000 ;
        878: q <= 32'b00000000000000000000000000000000 ;
        879: q <= 32'b00000000000000000000000000000000 ;
        880: q <= 32'b00000000000000000000000000000000 ;
        881: q <= 32'b00000000000000000000000000000000 ;
        882: q <= 32'b00000000000000000000000000000000 ;
        883: q <= 32'b00000000000000000000000000000000 ;
        884: q <= 32'b00000000000000000000000000000000 ;
        885: q <= 32'b00000000000000000000000000000000 ;
        886: q <= 32'b00000000000000000000000000000000 ;
        887: q <= 32'b00000000000000000000000000000000 ;
        888: q <= 32'b00000000000000000000000000000000 ;
        889: q <= 32'b00000000000000000000000000000000 ;
        890: q <= 32'b00000000000000000000000000000000 ;
        891: q <= 32'b00000000000000000000000000000000 ;
        892: q <= 32'b00000000000000000000000000000000 ;
        893: q <= 32'b00000000000000000000000000000000 ;
        894: q <= 32'b00000000000000000000000000000000 ;
        895: q <= 32'b00000000000000000000000000000000 ;
        896: q <= 32'b00000000000000000000000000000000 ;
        897: q <= 32'b00000000000000000000000000000000 ;
        898: q <= 32'b00000000000000000000000000000000 ;
        899: q <= 32'b00000000000000000000000000000000 ;
        900: q <= 32'b00000000000000000000000000000000 ;
        901: q <= 32'b00000000000000000000000000000000 ;
        902: q <= 32'b00000000000000000000000000000000 ;
        903: q <= 32'b00000000000000000000000000000000 ;
        904: q <= 32'b00000000000000000000000000000000 ;
        905: q <= 32'b00000000000000000000000000000000 ;
        906: q <= 32'b00000000000000000000000000000000 ;
        907: q <= 32'b00000000000000000000000000000000 ;
        908: q <= 32'b00000000000000000000000000000000 ;
        909: q <= 32'b00000000000000000000000000000000 ;
        910: q <= 32'b00000000000000000000000000000000 ;
        911: q <= 32'b00000000000000000000000000000000 ;
        912: q <= 32'b00000000000000000000000000000000 ;
        913: q <= 32'b00000000000000000000000000000000 ;
        914: q <= 32'b00000000000000000000000000000000 ;
        915: q <= 32'b00000000000000000000000000000000 ;
        916: q <= 32'b00000000000000000000000000000000 ;
        917: q <= 32'b00000000000000000000000000000000 ;
        918: q <= 32'b00000000000000000000000000000000 ;
        919: q <= 32'b00000000000000000000000000000000 ;
        920: q <= 32'b00000000000000000000000000000000 ;
        921: q <= 32'b00000000000000000000000000000000 ;
        922: q <= 32'b00000000000000000000000000000000 ;
        923: q <= 32'b00000000000000000000000000000000 ;
        924: q <= 32'b00000000000000000000000000000000 ;
        925: q <= 32'b00000000000000000000000000000000 ;
        926: q <= 32'b00000000000000000000000000000000 ;
        927: q <= 32'b00000000000000000000000000000000 ;
        928: q <= 32'b00000000000000000000000000000000 ;
        929: q <= 32'b00000000000000000000000000000000 ;
        930: q <= 32'b00000000000000000000000000000000 ;
        931: q <= 32'b00000000000000000000000000000000 ;
        932: q <= 32'b00000000000000000000000000000000 ;
        933: q <= 32'b00000000000000000000000000000000 ;
        934: q <= 32'b00000000000000000000000000000000 ;
        935: q <= 32'b00000000000000000000000000000000 ;
        936: q <= 32'b00000000000000000000000000000000 ;
        937: q <= 32'b00000000000000000000000000000000 ;
        938: q <= 32'b00000000000000000000000000000000 ;
        939: q <= 32'b00000000000000000000000000000000 ;
        940: q <= 32'b00000000000000000000000000000000 ;
        941: q <= 32'b00000000000000000000000000000000 ;
        942: q <= 32'b00000000000000000000000000000000 ;
        943: q <= 32'b00000000000000000000000000000000 ;
        944: q <= 32'b00000000000000000000000000000000 ;
        945: q <= 32'b00000000000000000000000000000000 ;
        946: q <= 32'b00000000000000000000000000000000 ;
        947: q <= 32'b00000000000000000000000000000000 ;
        948: q <= 32'b00000000000000000000000000000000 ;
        949: q <= 32'b00000000000000000000000000000000 ;
        950: q <= 32'b00000000000000000000000000000000 ;
        951: q <= 32'b00000000000000000000000000000000 ;
        952: q <= 32'b00000000000000000000000000000000 ;
        953: q <= 32'b00000000000000000000000000000000 ;
        954: q <= 32'b00000000000000000000000000000000 ;
        955: q <= 32'b00000000000000000000000000000000 ;
        956: q <= 32'b00000000000000000000000000000000 ;
        957: q <= 32'b00000000000000000000000000000000 ;
        958: q <= 32'b00000000000000000000000000000000 ;
        959: q <= 32'b00000000000000000000000000000000 ;
        960: q <= 32'b00000000000000000000000000000000 ;
        961: q <= 32'b00000000000000000000000000000000 ;
        962: q <= 32'b00000000000000000000000000000000 ;
        963: q <= 32'b00000000000000000000000000000000 ;
        964: q <= 32'b00000000000000000000000000000000 ;
        965: q <= 32'b00000000000000000000000000000000 ;
        966: q <= 32'b00000000000000000000000000000000 ;
        967: q <= 32'b00000000000000000000000000000000 ;
        968: q <= 32'b00000000000000000000000000000000 ;
        969: q <= 32'b00000000000000000000000000000000 ;
        970: q <= 32'b00000000000000000000000000000000 ;
        971: q <= 32'b00000000000000000000000000000000 ;
        972: q <= 32'b00000000000000000000000000000000 ;
        973: q <= 32'b00000000000000000000000000000000 ;
        974: q <= 32'b00000000000000000000000000000000 ;
        975: q <= 32'b00000000000000000000000000000000 ;
        976: q <= 32'b00000000000000000000000000000000 ;
        977: q <= 32'b00000000000000000000000000000000 ;
        978: q <= 32'b00000000000000000000000000000000 ;
        979: q <= 32'b00000000000000000000000000000000 ;
        980: q <= 32'b00000000000000000000000000000000 ;
        981: q <= 32'b00000000000000000000000000000000 ;
        982: q <= 32'b00000000000000000000000000000000 ;
        983: q <= 32'b00000000000000000000000000000000 ;
        984: q <= 32'b00000000000000000000000000000000 ;
        985: q <= 32'b00000000000000000000000000000000 ;
        986: q <= 32'b00000000000000000000000000000000 ;
        987: q <= 32'b00000000000000000000000000000000 ;
        988: q <= 32'b00000000000000000000000000000000 ;
        989: q <= 32'b00000000000000000000000000000000 ;
        990: q <= 32'b00000000000000000000000000000000 ;
        991: q <= 32'b00000000000000000000000000000000 ;
        992: q <= 32'b00000000000000000000000000000000 ;
        993: q <= 32'b00000000000000000000000000000000 ;
        994: q <= 32'b00000000000000000000000000000000 ;
        995: q <= 32'b00000000000000000000000000000000 ;
        996: q <= 32'b00000000000000000000000000000000 ;
        997: q <= 32'b00000000000000000000000000000000 ;
        998: q <= 32'b00000000000000000000000000000000 ;
        999: q <= 32'b00000000000000000000000000000000 ;
        1000: q <= 32'b00000000000000000000000000000000 ;
        1001: q <= 32'b00000000000000000000000000000000 ;
        1002: q <= 32'b00000000000000000000000000000000 ;
        1003: q <= 32'b00000000000000000000000000000000 ;
        1004: q <= 32'b00000000000000000000000000000000 ;
        1005: q <= 32'b00000000000000000000000000000000 ;
        1006: q <= 32'b00000000000000000000000000000000 ;
        1007: q <= 32'b00000000000000000000000000000000 ;
        1008: q <= 32'b00000000000000000000000000000000 ;
        1009: q <= 32'b00000000000000000000000000000000 ;
        1010: q <= 32'b00000000000000000000000000000000 ;
        1011: q <= 32'b00000000000000000000000000000000 ;
        1012: q <= 32'b00000000000000000000000000000000 ;
        1013: q <= 32'b00000000000000000000000000000000 ;
        1014: q <= 32'b00000000000000000000000000000000 ;
        1015: q <= 32'b00000000000000000000000000000000 ;
        1016: q <= 32'b00000000000000000000000000000000 ;
        1017: q <= 32'b00000000000000000000000000000000 ;
        1018: q <= 32'b00000000000000000000000000000000 ;
        1019: q <= 32'b00000000000000000000000000000000 ;
        1020: q <= 32'b00000000000000000000000000000000 ;
        1021: q <= 32'b00000000000000000000000000000000 ;
        1022: q <= 32'b00000000000000000000000000000000 ;
        1023: q <= 32'b00000000000000000000000000000000 ;
        default: q <= 32'b00000000000000000000000000000000;
    endcase
end

endmodule
