module mem_rom_weight_middle_01 (clock, address, q) ;
parameter DATA_WIDTH =  32;
input clock;
input [11:0] address;
output [DATA_WIDTH-1:0] q;
reg    [DATA_WIDTH-1:0] q;
always@(posedge clock) begin 
    case(address)
        0: q <= 32'b00111101100110000111101000000100 ;
        1: q <= 32'b00111101001100101111101010000110 ;
        2: q <= 32'b10111100100111010110010111000101 ;
        3: q <= 32'b00111100101111001010010010011001 ;
        4: q <= 32'b00111101110000111101101000101001 ;
        5: q <= 32'b00111011111010101111000110011110 ;
        6: q <= 32'b10111011000010111100110101111000 ;
        7: q <= 32'b00111101101101010011010101001110 ;
        8: q <= 32'b00111101101101001110011101110011 ;
        9: q <= 32'b00111101011011111111101011011100 ;
        10: q <= 32'b10111101100010001111101101010001 ;
        11: q <= 32'b00111101010101111010011100001101 ;
        12: q <= 32'b00111101010010111101110110001100 ;
        13: q <= 32'b10111100000001000100011101011011 ;
        14: q <= 32'b00111101101000001111110111010110 ;
        15: q <= 32'b00111101001011100011000110010000 ;
        16: q <= 32'b10111011101011100010110101110111 ;
        17: q <= 32'b00111100011110011101010000111110 ;
        18: q <= 32'b00111101011001011010010001111010 ;
        19: q <= 32'b00111101101110111001111111010010 ;
        20: q <= 32'b00111101100000101100011100101010 ;
        21: q <= 32'b10111101011111011101001111111011 ;
        22: q <= 32'b00111101100000001100111100010010 ;
        23: q <= 32'b00111101101000010100000111000011 ;
        24: q <= 32'b00111101100010011010110011000011 ;
        25: q <= 32'b00111101000110110010111101000000 ;
        26: q <= 32'b00111101101000011001000011000110 ;
        27: q <= 32'b10111101010110100111001001010011 ;
        28: q <= 32'b00111101110001011111001100110010 ;
        29: q <= 32'b10111101001110100001100001110101 ;
        30: q <= 32'b00111101100010000011101011101100 ;
        31: q <= 32'b10111100100110110101110000010100 ;
        32: q <= 32'b10111101101000001010100011100010 ;
        33: q <= 32'b10111101001011101011011001111111 ;
        34: q <= 32'b10111101101001011101111001100101 ;
        35: q <= 32'b00111101000100010111001111101111 ;
        36: q <= 32'b00111101110001011010111100101011 ;
        37: q <= 32'b10111101101101101111111101000011 ;
        38: q <= 32'b00111101001101001110000100111110 ;
        39: q <= 32'b10111011000111010110001110110100 ;
        40: q <= 32'b10111100101011100111101111000010 ;
        41: q <= 32'b00111011101011010010001000100000 ;
        42: q <= 32'b00111100011101010001101001010101 ;
        43: q <= 32'b00111100010001110000011001100010 ;
        44: q <= 32'b10111011000001110111110101100111 ;
        45: q <= 32'b10111101101001100111111011101000 ;
        46: q <= 32'b10111101001100110000011110000100 ;
        47: q <= 32'b00111101011001110011001000011000 ;
        48: q <= 32'b00111100111011010100001010100001 ;
        49: q <= 32'b00111101110000010001010100011001 ;
        50: q <= 32'b10111101110010111011100110100100 ;
        51: q <= 32'b00111101101101101010111010110010 ;
        52: q <= 32'b00111101110110100110000011000000 ;
        53: q <= 32'b10111101000100110010111010000010 ;
        54: q <= 32'b00111101010101001100101101111110 ;
        55: q <= 32'b10111101010001111001110111110000 ;
        56: q <= 32'b00111100100010101010010110110000 ;
        57: q <= 32'b10111101100000111000001110111001 ;
        58: q <= 32'b00111101101010011110001100001100 ;
        59: q <= 32'b00111001100010000001001101100111 ;
        60: q <= 32'b00111100110110100111110001000101 ;
        61: q <= 32'b10111100100001100011110100111001 ;
        62: q <= 32'b00111101100011011011100101000000 ;
        63: q <= 32'b00111101100100001010011111010000 ;
        64: q <= 32'b00111101100011000100010001111010 ;
        65: q <= 32'b10111100001101111001100111100111 ;
        66: q <= 32'b10111010110111100101100100100110 ;
        67: q <= 32'b10111101001100000001101110010000 ;
        68: q <= 32'b10111101000100101100000011100011 ;
        69: q <= 32'b10111100110111100010001101101001 ;
        70: q <= 32'b00111100000011010010010011101100 ;
        71: q <= 32'b10111101100110001011001110010100 ;
        72: q <= 32'b00111101000111010000100101100000 ;
        73: q <= 32'b10111101100100110100101110010110 ;
        74: q <= 32'b00111101100001011100100110110011 ;
        75: q <= 32'b10111010111111011011010011010010 ;
        76: q <= 32'b10111100111101010101100110100101 ;
        77: q <= 32'b10111101101100101110001110000100 ;
        78: q <= 32'b00111110000000000001001011110111 ;
        79: q <= 32'b10111100110101111010100100011010 ;
        80: q <= 32'b00111011111101100101110110110101 ;
        81: q <= 32'b00111101011101000101100110110011 ;
        82: q <= 32'b00111101101010001111000011000001 ;
        83: q <= 32'b00111101111000010101000110000011 ;
        84: q <= 32'b00111100001110100110011011011010 ;
        85: q <= 32'b10111101100111011101001101110101 ;
        86: q <= 32'b00111101011100001101011110010110 ;
        87: q <= 32'b00111100111111000110110110001000 ;
        88: q <= 32'b10111100100001000111011010110111 ;
        89: q <= 32'b00111101100011101111110110000100 ;
        90: q <= 32'b10111101100000011111101101101110 ;
        91: q <= 32'b10111101011100011100010101001100 ;
        92: q <= 32'b00111101100101110110011111010010 ;
        93: q <= 32'b00111100100110000101110000011100 ;
        94: q <= 32'b00111100011111110110010110111111 ;
        95: q <= 32'b00111011100011101100010100011100 ;
        96: q <= 32'b00111100101110110101110111000111 ;
        97: q <= 32'b10111100011110001111001110000001 ;
        98: q <= 32'b10111101100001101000101011011111 ;
        99: q <= 32'b10111101100000001110001101110111 ;
        100: q <= 32'b10111100101011010111000001001111 ;
        101: q <= 32'b00111100010110000001101001111110 ;
        102: q <= 32'b10111101000111100101001001011111 ;
        103: q <= 32'b00111101101110000000110111000010 ;
        104: q <= 32'b00000000000000000000000000000000 ;
        105: q <= 32'b00000000000000000000000000000000 ;
        106: q <= 32'b00000000000000000000000000000000 ;
        107: q <= 32'b00000000000000000000000000000000 ;
        108: q <= 32'b00000000000000000000000000000000 ;
        109: q <= 32'b00000000000000000000000000000000 ;
        110: q <= 32'b00000000000000000000000000000000 ;
        111: q <= 32'b00000000000000000000000000000000 ;
        112: q <= 32'b00000000000000000000000000000000 ;
        113: q <= 32'b00000000000000000000000000000000 ;
        114: q <= 32'b00000000000000000000000000000000 ;
        115: q <= 32'b00000000000000000000000000000000 ;
        116: q <= 32'b00000000000000000000000000000000 ;
        117: q <= 32'b00000000000000000000000000000000 ;
        118: q <= 32'b00000000000000000000000000000000 ;
        119: q <= 32'b00000000000000000000000000000000 ;
        120: q <= 32'b00000000000000000000000000000000 ;
        121: q <= 32'b00000000000000000000000000000000 ;
        122: q <= 32'b00000000000000000000000000000000 ;
        123: q <= 32'b00000000000000000000000000000000 ;
        124: q <= 32'b00000000000000000000000000000000 ;
        125: q <= 32'b00000000000000000000000000000000 ;
        126: q <= 32'b00000000000000000000000000000000 ;
        127: q <= 32'b00000000000000000000000000000000 ;
        128: q <= 32'b00111100110101000101110001110011 ;
        129: q <= 32'b00111101010111011010111111010101 ;
        130: q <= 32'b10111101100001111100010110010011 ;
        131: q <= 32'b00111110010000100010001100011000 ;
        132: q <= 32'b00111100101101001100111100111111 ;
        133: q <= 32'b10111101000101000011111001011011 ;
        134: q <= 32'b10111101100111000101000111110011 ;
        135: q <= 32'b10111101000010000100000011111111 ;
        136: q <= 32'b00111101001001011011011111001000 ;
        137: q <= 32'b00111100011000000010111110010001 ;
        138: q <= 32'b00111101000001100000111011010011 ;
        139: q <= 32'b00111101001101011101000100000010 ;
        140: q <= 32'b00111101001101111101001111100111 ;
        141: q <= 32'b10111101100001011111100001111001 ;
        142: q <= 32'b10111101100011010100100001100110 ;
        143: q <= 32'b10111101001000110010101001000110 ;
        144: q <= 32'b10111101010001111001110001011010 ;
        145: q <= 32'b00111101000011000100101110001010 ;
        146: q <= 32'b10111101111100011101011001011101 ;
        147: q <= 32'b00111110000100100000111101100001 ;
        148: q <= 32'b00111101011100110001110111000011 ;
        149: q <= 32'b00111100111010100110011011000101 ;
        150: q <= 32'b10111101001100110001001001001011 ;
        151: q <= 32'b10111110001100100010110100001110 ;
        152: q <= 32'b10111101011110101110001000000111 ;
        153: q <= 32'b00111101000100011100011101001110 ;
        154: q <= 32'b10111101000100001000110101010111 ;
        155: q <= 32'b00111101001101000001001001000111 ;
        156: q <= 32'b10111101111100101001010100010000 ;
        157: q <= 32'b10111100011010101100010000111101 ;
        158: q <= 32'b10111101100010011111000101111111 ;
        159: q <= 32'b10111101110001110001000110000101 ;
        160: q <= 32'b00111101100110001111011111100000 ;
        161: q <= 32'b00111100111100111010011000101000 ;
        162: q <= 32'b00111101100111001010010001001000 ;
        163: q <= 32'b10111101001100100110000101011100 ;
        164: q <= 32'b00111100111001010111001101011001 ;
        165: q <= 32'b00111101011000110111101011101100 ;
        166: q <= 32'b10111101101010101101001100110100 ;
        167: q <= 32'b10111101100110001101111101011101 ;
        168: q <= 32'b10111101111110100000010111000001 ;
        169: q <= 32'b10111100000001111011100000010101 ;
        170: q <= 32'b10111110000100110111100100111010 ;
        171: q <= 32'b00111101001111111110010010100000 ;
        172: q <= 32'b00111101101000110010010010001111 ;
        173: q <= 32'b10111100011110111110010011010000 ;
        174: q <= 32'b00111011101110000011100000100011 ;
        175: q <= 32'b10111101101010000101001111011011 ;
        176: q <= 32'b00111100100010010100111100101101 ;
        177: q <= 32'b00111101110110010001001010001110 ;
        178: q <= 32'b10111101001010101011001110110000 ;
        179: q <= 32'b10111100100101001110101010001010 ;
        180: q <= 32'b10111101011111010010011111111101 ;
        181: q <= 32'b10111101001011100000010010111101 ;
        182: q <= 32'b10111101011110011000010001001010 ;
        183: q <= 32'b10111101100000010010000110001111 ;
        184: q <= 32'b00111101000100011000100000111001 ;
        185: q <= 32'b10111100101011001111000011111100 ;
        186: q <= 32'b10111011000011101011010001110101 ;
        187: q <= 32'b10111101101001000010101100101010 ;
        188: q <= 32'b10111101010000000110000110110111 ;
        189: q <= 32'b10111101100101100100001010011011 ;
        190: q <= 32'b00111101100100101100100110001010 ;
        191: q <= 32'b00111101101011101000001111111011 ;
        192: q <= 32'b00111101111000010011101101111011 ;
        193: q <= 32'b10111101101111010000101010010010 ;
        194: q <= 32'b10111101111110000000111111100111 ;
        195: q <= 32'b00111101011010001111111101110101 ;
        196: q <= 32'b10111101010111000000111111101000 ;
        197: q <= 32'b00111101001000001011101110011110 ;
        198: q <= 32'b00111100011110011111110111110000 ;
        199: q <= 32'b10111101001101011010110111101011 ;
        200: q <= 32'b10111101011001110010001010000110 ;
        201: q <= 32'b00111101001110000100000101100110 ;
        202: q <= 32'b00111100011011111111000001100010 ;
        203: q <= 32'b10111101100110111100101000010001 ;
        204: q <= 32'b00111101011010010101111111111111 ;
        205: q <= 32'b10111101100110011000001111101111 ;
        206: q <= 32'b10111100101111111001111000101000 ;
        207: q <= 32'b10111110011000100001011000100101 ;
        208: q <= 32'b00111110010001000101100110101111 ;
        209: q <= 32'b10111100100110110010000100001101 ;
        210: q <= 32'b10111101100000011111001010011010 ;
        211: q <= 32'b00111101101001111110000101011001 ;
        212: q <= 32'b00111101000110110101001001111001 ;
        213: q <= 32'b10111101111000001101100010001001 ;
        214: q <= 32'b00111101101010010110110010101111 ;
        215: q <= 32'b00111101000100110011100101001001 ;
        216: q <= 32'b10111100110011101011100000011101 ;
        217: q <= 32'b10111101011010001001110110000101 ;
        218: q <= 32'b10111101010101010000110000111010 ;
        219: q <= 32'b10111101101100010000100110010011 ;
        220: q <= 32'b10111101010000011011100001100100 ;
        221: q <= 32'b00111101100101111111001011001000 ;
        222: q <= 32'b00111101000000111010111001111000 ;
        223: q <= 32'b00111101100111010000010111111100 ;
        224: q <= 32'b10111100000101001111001010111000 ;
        225: q <= 32'b10111101010011011100011110111001 ;
        226: q <= 32'b10111101011010011011011001001001 ;
        227: q <= 32'b00111101011111111011011000111111 ;
        228: q <= 32'b10111101101011110110011111111111 ;
        229: q <= 32'b00111101010000110000011101100110 ;
        230: q <= 32'b00111101101111101000001111101001 ;
        231: q <= 32'b00111101100111101110101110111110 ;
        232: q <= 32'b00000000000000000000000000000000 ;
        233: q <= 32'b00000000000000000000000000000000 ;
        234: q <= 32'b00000000000000000000000000000000 ;
        235: q <= 32'b00000000000000000000000000000000 ;
        236: q <= 32'b00000000000000000000000000000000 ;
        237: q <= 32'b00000000000000000000000000000000 ;
        238: q <= 32'b00000000000000000000000000000000 ;
        239: q <= 32'b00000000000000000000000000000000 ;
        240: q <= 32'b00000000000000000000000000000000 ;
        241: q <= 32'b00000000000000000000000000000000 ;
        242: q <= 32'b00000000000000000000000000000000 ;
        243: q <= 32'b00000000000000000000000000000000 ;
        244: q <= 32'b00000000000000000000000000000000 ;
        245: q <= 32'b00000000000000000000000000000000 ;
        246: q <= 32'b00000000000000000000000000000000 ;
        247: q <= 32'b00000000000000000000000000000000 ;
        248: q <= 32'b00000000000000000000000000000000 ;
        249: q <= 32'b00000000000000000000000000000000 ;
        250: q <= 32'b00000000000000000000000000000000 ;
        251: q <= 32'b00000000000000000000000000000000 ;
        252: q <= 32'b00000000000000000000000000000000 ;
        253: q <= 32'b00000000000000000000000000000000 ;
        254: q <= 32'b00000000000000000000000000000000 ;
        255: q <= 32'b00000000000000000000000000000000 ;
        256: q <= 32'b00111101010011100000100101101110 ;
        257: q <= 32'b00111101110001001000101010100101 ;
        258: q <= 32'b00111100010001111111110100100101 ;
        259: q <= 32'b10111101001011111111011101000011 ;
        260: q <= 32'b10111110000011010011110011111011 ;
        261: q <= 32'b10111101001001001111010011000001 ;
        262: q <= 32'b00111110001011010101100110101101 ;
        263: q <= 32'b10111101110010000100111001000110 ;
        264: q <= 32'b10111101101111101111101101101011 ;
        265: q <= 32'b00111100011111110110001001101101 ;
        266: q <= 32'b10111101100111111111100100000001 ;
        267: q <= 32'b00111100001111101100110110000100 ;
        268: q <= 32'b10111100100001000101011000010100 ;
        269: q <= 32'b00111101000000100000011001010110 ;
        270: q <= 32'b00111100100001000000111001001111 ;
        271: q <= 32'b10111101110110101100101101111001 ;
        272: q <= 32'b00111110000001111100000100111100 ;
        273: q <= 32'b00111101111100001001000110101110 ;
        274: q <= 32'b00111101000010110001010101101101 ;
        275: q <= 32'b10111110010000100100110000110001 ;
        276: q <= 32'b00111011001110010110001100000001 ;
        277: q <= 32'b10111101010011001100100011010010 ;
        278: q <= 32'b10111100110110100001000100101011 ;
        279: q <= 32'b10111011110010000000110010010010 ;
        280: q <= 32'b00111110000010100000000101101101 ;
        281: q <= 32'b00111010111101110001100101011110 ;
        282: q <= 32'b00111100110001101000100111100000 ;
        283: q <= 32'b10111101000011100011111000001001 ;
        284: q <= 32'b10111100101010011001100111100000 ;
        285: q <= 32'b00111011110101100110001111011101 ;
        286: q <= 32'b00111100111100001101010011100000 ;
        287: q <= 32'b00111101010111011101111001110100 ;
        288: q <= 32'b10111101000100111000011101101000 ;
        289: q <= 32'b10111101100011101110010001111011 ;
        290: q <= 32'b10111100110101010010010000101101 ;
        291: q <= 32'b10111100101111110011010100100011 ;
        292: q <= 32'b10111101001100100100010111011011 ;
        293: q <= 32'b00111101101000011111011100011100 ;
        294: q <= 32'b10111100110101111101010101011011 ;
        295: q <= 32'b00111100001110100111101101100010 ;
        296: q <= 32'b10111011111001110111110001100011 ;
        297: q <= 32'b10111100011101001000100000110110 ;
        298: q <= 32'b00111101100011101011001110101100 ;
        299: q <= 32'b00111110000000110001110101111011 ;
        300: q <= 32'b00111101000000010111000011110100 ;
        301: q <= 32'b10111101110101000011110111001010 ;
        302: q <= 32'b10111100100010101111001100101011 ;
        303: q <= 32'b00111101100101100110011111111110 ;
        304: q <= 32'b00111011000010110101001011100010 ;
        305: q <= 32'b10111101111011100111111100101111 ;
        306: q <= 32'b00111100111010011100010000001011 ;
        307: q <= 32'b00111100011011000001100101110000 ;
        308: q <= 32'b10111101100000010010101010010010 ;
        309: q <= 32'b00111001111111011000011001010010 ;
        310: q <= 32'b00111101100111101111001010101000 ;
        311: q <= 32'b00111101101011011100110011001101 ;
        312: q <= 32'b10111101000000100001011011011000 ;
        313: q <= 32'b10111101010000001000100100110101 ;
        314: q <= 32'b10111101100001100001110001110110 ;
        315: q <= 32'b00111101100100100110010111001011 ;
        316: q <= 32'b10111101110010011101110101101100 ;
        317: q <= 32'b10111001001100110111010001110110 ;
        318: q <= 32'b10111110000110101101000010001000 ;
        319: q <= 32'b00111110000011110010001000011101 ;
        320: q <= 32'b10111100101111101101011010001010 ;
        321: q <= 32'b00111011011101110100000100101101 ;
        322: q <= 32'b00111101101000011100110000001110 ;
        323: q <= 32'b00111100100000011001101010101000 ;
        324: q <= 32'b10111101000111100111010001001001 ;
        325: q <= 32'b00111100111100100010001011011010 ;
        326: q <= 32'b00111100101101000010101011110011 ;
        327: q <= 32'b10111101100011101010100101100001 ;
        328: q <= 32'b00111010000100010010000110111011 ;
        329: q <= 32'b00111101110111000001110101100000 ;
        330: q <= 32'b00111100101100010001000101101111 ;
        331: q <= 32'b10111010001101111001100101001100 ;
        332: q <= 32'b00111101100010110111100101101001 ;
        333: q <= 32'b00111101001110100001110011011000 ;
        334: q <= 32'b10111100011011101010010000011101 ;
        335: q <= 32'b00111101101100010111010000110010 ;
        336: q <= 32'b00111011000000101100110001100011 ;
        337: q <= 32'b00111101101111010100010000100000 ;
        338: q <= 32'b00111011101110010101000110111000 ;
        339: q <= 32'b00111101111001100100110000001111 ;
        340: q <= 32'b00111101111110101011001000001111 ;
        341: q <= 32'b10111101100110011001001100000010 ;
        342: q <= 32'b10111100011110101101010010100001 ;
        343: q <= 32'b10111101010110111011110110001000 ;
        344: q <= 32'b00111100110001000111111011101110 ;
        345: q <= 32'b00111101100110111101011011100000 ;
        346: q <= 32'b00111101101101110111111101110011 ;
        347: q <= 32'b10111100100011110111010010101111 ;
        348: q <= 32'b10111100010111111001111000111101 ;
        349: q <= 32'b00111011010111011111011011011101 ;
        350: q <= 32'b10111011101001010001101100101000 ;
        351: q <= 32'b00111101010001111101010110111000 ;
        352: q <= 32'b00111101100100011101101110001011 ;
        353: q <= 32'b00111101000001000010110010011101 ;
        354: q <= 32'b00111101100110101110101100001010 ;
        355: q <= 32'b00111110001110111001010100001101 ;
        356: q <= 32'b10111010100111010010011000010100 ;
        357: q <= 32'b10111011100100011010110001000001 ;
        358: q <= 32'b00111101001001000101110111001010 ;
        359: q <= 32'b00111101101100011010001111010010 ;
        360: q <= 32'b00000000000000000000000000000000 ;
        361: q <= 32'b00000000000000000000000000000000 ;
        362: q <= 32'b00000000000000000000000000000000 ;
        363: q <= 32'b00000000000000000000000000000000 ;
        364: q <= 32'b00000000000000000000000000000000 ;
        365: q <= 32'b00000000000000000000000000000000 ;
        366: q <= 32'b00000000000000000000000000000000 ;
        367: q <= 32'b00000000000000000000000000000000 ;
        368: q <= 32'b00000000000000000000000000000000 ;
        369: q <= 32'b00000000000000000000000000000000 ;
        370: q <= 32'b00000000000000000000000000000000 ;
        371: q <= 32'b00000000000000000000000000000000 ;
        372: q <= 32'b00000000000000000000000000000000 ;
        373: q <= 32'b00000000000000000000000000000000 ;
        374: q <= 32'b00000000000000000000000000000000 ;
        375: q <= 32'b00000000000000000000000000000000 ;
        376: q <= 32'b00000000000000000000000000000000 ;
        377: q <= 32'b00000000000000000000000000000000 ;
        378: q <= 32'b00000000000000000000000000000000 ;
        379: q <= 32'b00000000000000000000000000000000 ;
        380: q <= 32'b00000000000000000000000000000000 ;
        381: q <= 32'b00000000000000000000000000000000 ;
        382: q <= 32'b00000000000000000000000000000000 ;
        383: q <= 32'b00000000000000000000000000000000 ;
        384: q <= 32'b00111101010001000110101111010010 ;
        385: q <= 32'b00111101100111111110110111000010 ;
        386: q <= 32'b10111110000010011111010101010001 ;
        387: q <= 32'b10111101100000111000001001101100 ;
        388: q <= 32'b10111101110101100111100000000000 ;
        389: q <= 32'b00111101001100111110001111110101 ;
        390: q <= 32'b10111101011010101101000101001001 ;
        391: q <= 32'b10111101000100111110000110100100 ;
        392: q <= 32'b10111101110110001110101001011100 ;
        393: q <= 32'b10111101001101101111100000011001 ;
        394: q <= 32'b00111100110110001011011101111010 ;
        395: q <= 32'b00111101101011000101111100110010 ;
        396: q <= 32'b10111101011111111110110101101000 ;
        397: q <= 32'b10111100100111111101100101010000 ;
        398: q <= 32'b00111100000110101000111111100011 ;
        399: q <= 32'b10111101100111011110001111101010 ;
        400: q <= 32'b00111100011100101000001001001101 ;
        401: q <= 32'b00111101111010010000000001010011 ;
        402: q <= 32'b10111101101011011111011001111110 ;
        403: q <= 32'b00111100100110000111111110111110 ;
        404: q <= 32'b00111100011111001000100001110101 ;
        405: q <= 32'b00111101111111011110001011111110 ;
        406: q <= 32'b10111100101001101111101001111000 ;
        407: q <= 32'b10111101101101001010011101011110 ;
        408: q <= 32'b10111101101011000000010100110100 ;
        409: q <= 32'b10111101100111000111001100111101 ;
        410: q <= 32'b10111101000001001001101011111000 ;
        411: q <= 32'b10111100111000000001010100011011 ;
        412: q <= 32'b10111110001000111101100001101010 ;
        413: q <= 32'b00111101100111001111011101011111 ;
        414: q <= 32'b10111101000101000010011100111001 ;
        415: q <= 32'b00111100100111101101100010010001 ;
        416: q <= 32'b10111101111010101000110010011101 ;
        417: q <= 32'b00111100100101100000111100101101 ;
        418: q <= 32'b00111101011010110011111110110111 ;
        419: q <= 32'b00111101110100110000110101111011 ;
        420: q <= 32'b10111101100111101010101000010111 ;
        421: q <= 32'b00111101100111010100011101101110 ;
        422: q <= 32'b10111100110100011011110100000011 ;
        423: q <= 32'b00111101101011011010000100010011 ;
        424: q <= 32'b00111101011101000110100011010101 ;
        425: q <= 32'b00111100111010011111111001001001 ;
        426: q <= 32'b00111101110111111101111100111011 ;
        427: q <= 32'b00111110001100110000001100000011 ;
        428: q <= 32'b10111110000000000001001100111011 ;
        429: q <= 32'b10111101101100011101101011010111 ;
        430: q <= 32'b00111101110000011110110111100010 ;
        431: q <= 32'b10111110000000111000101101111001 ;
        432: q <= 32'b10111100100010001001010101000000 ;
        433: q <= 32'b00111101011111101001000010001000 ;
        434: q <= 32'b00111101000111001011100101101001 ;
        435: q <= 32'b00111011011001111100011111110110 ;
        436: q <= 32'b10111100101110000110101111011110 ;
        437: q <= 32'b10111101001100100110011001011001 ;
        438: q <= 32'b10111110011100001000101111001110 ;
        439: q <= 32'b00111101101001000101001011000000 ;
        440: q <= 32'b10111101000100000111001011000110 ;
        441: q <= 32'b00111101000011101101001010100001 ;
        442: q <= 32'b10111100101101000011011011010101 ;
        443: q <= 32'b10111100100000100000101010101110 ;
        444: q <= 32'b10111101111010101101001101010000 ;
        445: q <= 32'b00111010010001100100011000001011 ;
        446: q <= 32'b10111100001111110110011001011100 ;
        447: q <= 32'b10111100000011101110011001111011 ;
        448: q <= 32'b00111101110010111101111001000100 ;
        449: q <= 32'b10111100100010100111000101001101 ;
        450: q <= 32'b10111110000100010101101100001110 ;
        451: q <= 32'b00111100100010110011101001001100 ;
        452: q <= 32'b00111011111010101001010011000101 ;
        453: q <= 32'b10111100010101010111111110010100 ;
        454: q <= 32'b00111101101111110000111110110010 ;
        455: q <= 32'b10111110000000000111101100010111 ;
        456: q <= 32'b00111101000010110010100001100001 ;
        457: q <= 32'b00111101011101011111100101100001 ;
        458: q <= 32'b00111100110110011100001000101111 ;
        459: q <= 32'b00111010100111100110000101111101 ;
        460: q <= 32'b00111101100100111001011101000101 ;
        461: q <= 32'b10111101011010110001011010111010 ;
        462: q <= 32'b00111110000010010010011101000001 ;
        463: q <= 32'b10111101101110011110101001101000 ;
        464: q <= 32'b10111101000011100111111010110100 ;
        465: q <= 32'b10111101001100110111010101010000 ;
        466: q <= 32'b00111110000100111010001000010101 ;
        467: q <= 32'b10111100111001000101000111011001 ;
        468: q <= 32'b10111110001011010100001100000111 ;
        469: q <= 32'b10111101000001111111101100110001 ;
        470: q <= 32'b10111101000000111111101100010101 ;
        471: q <= 32'b10111101010010011100100110011001 ;
        472: q <= 32'b00111100101100000011110011110100 ;
        473: q <= 32'b10111011111101000110101101100100 ;
        474: q <= 32'b00111101000010001100010100110100 ;
        475: q <= 32'b10111101100000010010100100101011 ;
        476: q <= 32'b10111101011011101001110100010011 ;
        477: q <= 32'b00111110000111111101010110101111 ;
        478: q <= 32'b00111101100110101011000011110101 ;
        479: q <= 32'b00111101010001110011111100011011 ;
        480: q <= 32'b00111101001001111001110010000001 ;
        481: q <= 32'b10111101010000100100100101001011 ;
        482: q <= 32'b10111101000010000010111001001111 ;
        483: q <= 32'b00111101100010010000010100110000 ;
        484: q <= 32'b10111101110001101010010111011100 ;
        485: q <= 32'b00111110000001101101111110101001 ;
        486: q <= 32'b00111101100110110101100110011101 ;
        487: q <= 32'b00111101101010000001000010101011 ;
        488: q <= 32'b00000000000000000000000000000000 ;
        489: q <= 32'b00000000000000000000000000000000 ;
        490: q <= 32'b00000000000000000000000000000000 ;
        491: q <= 32'b00000000000000000000000000000000 ;
        492: q <= 32'b00000000000000000000000000000000 ;
        493: q <= 32'b00000000000000000000000000000000 ;
        494: q <= 32'b00000000000000000000000000000000 ;
        495: q <= 32'b00000000000000000000000000000000 ;
        496: q <= 32'b00000000000000000000000000000000 ;
        497: q <= 32'b00000000000000000000000000000000 ;
        498: q <= 32'b00000000000000000000000000000000 ;
        499: q <= 32'b00000000000000000000000000000000 ;
        500: q <= 32'b00000000000000000000000000000000 ;
        501: q <= 32'b00000000000000000000000000000000 ;
        502: q <= 32'b00000000000000000000000000000000 ;
        503: q <= 32'b00000000000000000000000000000000 ;
        504: q <= 32'b00000000000000000000000000000000 ;
        505: q <= 32'b00000000000000000000000000000000 ;
        506: q <= 32'b00000000000000000000000000000000 ;
        507: q <= 32'b00000000000000000000000000000000 ;
        508: q <= 32'b00000000000000000000000000000000 ;
        509: q <= 32'b00000000000000000000000000000000 ;
        510: q <= 32'b00000000000000000000000000000000 ;
        511: q <= 32'b00000000000000000000000000000000 ;
        512: q <= 32'b00111101010110001111101011100111 ;
        513: q <= 32'b00111011010011100110100101100110 ;
        514: q <= 32'b10111101000000001101010011111001 ;
        515: q <= 32'b00111110000001111000010011011010 ;
        516: q <= 32'b00111101101011110000001100100100 ;
        517: q <= 32'b10111101111110101001100110110011 ;
        518: q <= 32'b10111100100111100011101100101010 ;
        519: q <= 32'b10111100000110000101101110011010 ;
        520: q <= 32'b10111101110011010000100000000110 ;
        521: q <= 32'b10111101101011011110001111001100 ;
        522: q <= 32'b10111101001011110100000001011110 ;
        523: q <= 32'b00111101100101001000111011110001 ;
        524: q <= 32'b10111100110100110111001000000010 ;
        525: q <= 32'b00111100110101000010110111001100 ;
        526: q <= 32'b10111100001101010011000011101010 ;
        527: q <= 32'b00111101101101101011010111000001 ;
        528: q <= 32'b00111101010001110010110100011010 ;
        529: q <= 32'b00111100100111100000100001011111 ;
        530: q <= 32'b00111101000101100111000110011110 ;
        531: q <= 32'b00111101110100011110100010001100 ;
        532: q <= 32'b10111101110000110100100101101011 ;
        533: q <= 32'b00111100001001101011111101110010 ;
        534: q <= 32'b00111100001011100100010100101100 ;
        535: q <= 32'b10111100111111011000001010010111 ;
        536: q <= 32'b10111101110101101101010111111000 ;
        537: q <= 32'b10111101011011111100001110011100 ;
        538: q <= 32'b00111101101110011001010110001011 ;
        539: q <= 32'b00111101101001100000000111001100 ;
        540: q <= 32'b00111100100100001010001100100000 ;
        541: q <= 32'b00111110010000011100100010110100 ;
        542: q <= 32'b00111101000111101101010000110110 ;
        543: q <= 32'b10111101001010000101010011001010 ;
        544: q <= 32'b00111101011001101100011111111100 ;
        545: q <= 32'b10111101100110101111100101100111 ;
        546: q <= 32'b00111011000001110000111101101101 ;
        547: q <= 32'b10111100001111111101011110111100 ;
        548: q <= 32'b10111101001110101011100010101111 ;
        549: q <= 32'b10111101011011001000000000111111 ;
        550: q <= 32'b10111101110111101100001011011010 ;
        551: q <= 32'b00111101011001001111010011101110 ;
        552: q <= 32'b10111101111011010000110000100011 ;
        553: q <= 32'b00111101100101111101001001101110 ;
        554: q <= 32'b10111101101101101110000011100100 ;
        555: q <= 32'b10111100100010001110110001010111 ;
        556: q <= 32'b10111100110111100100010011100000 ;
        557: q <= 32'b00111101100101110110110011011001 ;
        558: q <= 32'b10111101100010000111000000000011 ;
        559: q <= 32'b00111010000001100000101010110111 ;
        560: q <= 32'b10111100110010011100001000101000 ;
        561: q <= 32'b00111100010010000010010011100100 ;
        562: q <= 32'b10111101101000011110100100011001 ;
        563: q <= 32'b00111101011101011010111001011001 ;
        564: q <= 32'b10111101010011100001111011010000 ;
        565: q <= 32'b00111101000001110101100101001010 ;
        566: q <= 32'b00111011010110111011100101011000 ;
        567: q <= 32'b00111110001100100001101110111111 ;
        568: q <= 32'b10111101000111000100000110100000 ;
        569: q <= 32'b10111101001000001100111011010000 ;
        570: q <= 32'b10111101010101010011011011000011 ;
        571: q <= 32'b00111101001100111000010110010011 ;
        572: q <= 32'b00111101001101111100010100010100 ;
        573: q <= 32'b00111101001011110110111011111101 ;
        574: q <= 32'b10111100101110000110011101111111 ;
        575: q <= 32'b00111101101011010100101100001001 ;
        576: q <= 32'b00111100001110110100010001010101 ;
        577: q <= 32'b10111100011001001011010011011100 ;
        578: q <= 32'b10111101010110011111101000110010 ;
        579: q <= 32'b00111100111101101111111100011100 ;
        580: q <= 32'b10111101110010010000000110000111 ;
        581: q <= 32'b00111101110001010101111000111101 ;
        582: q <= 32'b00111011110111011010010011100111 ;
        583: q <= 32'b10111100001100001111011010010111 ;
        584: q <= 32'b00111101010001010110110011010101 ;
        585: q <= 32'b10111100111001101101001110100011 ;
        586: q <= 32'b10111101000111000101110011010010 ;
        587: q <= 32'b00111010011101110010100100100001 ;
        588: q <= 32'b00111101000000010001011100110110 ;
        589: q <= 32'b00111100110000101100111001000010 ;
        590: q <= 32'b00111101001000110000001101110001 ;
        591: q <= 32'b10111101111100001001001011101001 ;
        592: q <= 32'b00111101110111001001100100100111 ;
        593: q <= 32'b00111110000101000010010010100111 ;
        594: q <= 32'b10111101110010100101001011111101 ;
        595: q <= 32'b00111101001101010011010100001001 ;
        596: q <= 32'b00111101101010111010111101000110 ;
        597: q <= 32'b00111011000101110101011111101011 ;
        598: q <= 32'b00111100101001110111101010000000 ;
        599: q <= 32'b10111101011001100111011001110100 ;
        600: q <= 32'b10111101011000110000000111011000 ;
        601: q <= 32'b10111100111010110010000010100000 ;
        602: q <= 32'b00111101101011110100011001011101 ;
        603: q <= 32'b00111101100010011100010100001010 ;
        604: q <= 32'b10111101010111100101101001101011 ;
        605: q <= 32'b10111100111111100001011111110001 ;
        606: q <= 32'b00111101000100000001011010010011 ;
        607: q <= 32'b00111101100000000000100000000110 ;
        608: q <= 32'b00111101010101011001101110101101 ;
        609: q <= 32'b00111100000101101001111100011111 ;
        610: q <= 32'b00111100110110000000010000001111 ;
        611: q <= 32'b00111101011000111000001001011111 ;
        612: q <= 32'b00111000101001101011011000001110 ;
        613: q <= 32'b10111101101100001010000000100101 ;
        614: q <= 32'b00111011101010111111001110011100 ;
        615: q <= 32'b10111101011010111111101000000100 ;
        616: q <= 32'b00000000000000000000000000000000 ;
        617: q <= 32'b00000000000000000000000000000000 ;
        618: q <= 32'b00000000000000000000000000000000 ;
        619: q <= 32'b00000000000000000000000000000000 ;
        620: q <= 32'b00000000000000000000000000000000 ;
        621: q <= 32'b00000000000000000000000000000000 ;
        622: q <= 32'b00000000000000000000000000000000 ;
        623: q <= 32'b00000000000000000000000000000000 ;
        624: q <= 32'b00000000000000000000000000000000 ;
        625: q <= 32'b00000000000000000000000000000000 ;
        626: q <= 32'b00000000000000000000000000000000 ;
        627: q <= 32'b00000000000000000000000000000000 ;
        628: q <= 32'b00000000000000000000000000000000 ;
        629: q <= 32'b00000000000000000000000000000000 ;
        630: q <= 32'b00000000000000000000000000000000 ;
        631: q <= 32'b00000000000000000000000000000000 ;
        632: q <= 32'b00000000000000000000000000000000 ;
        633: q <= 32'b00000000000000000000000000000000 ;
        634: q <= 32'b00000000000000000000000000000000 ;
        635: q <= 32'b00000000000000000000000000000000 ;
        636: q <= 32'b00000000000000000000000000000000 ;
        637: q <= 32'b00000000000000000000000000000000 ;
        638: q <= 32'b00000000000000000000000000000000 ;
        639: q <= 32'b00000000000000000000000000000000 ;
        640: q <= 32'b00111010001011010011101100011001 ;
        641: q <= 32'b10111110001001111011101001001011 ;
        642: q <= 32'b10111011010010100101010001111101 ;
        643: q <= 32'b00111101100011010100010100110111 ;
        644: q <= 32'b00111101110010000111100010011011 ;
        645: q <= 32'b00111100101000000000001001000100 ;
        646: q <= 32'b00111101101111100100111010100111 ;
        647: q <= 32'b00111101100101001010010011100000 ;
        648: q <= 32'b10111101110000000001001110011101 ;
        649: q <= 32'b00111011011100000100101100100001 ;
        650: q <= 32'b10111100101110010010011001000001 ;
        651: q <= 32'b10111101100111100101011001001110 ;
        652: q <= 32'b00111101100100110010000011011100 ;
        653: q <= 32'b10111101111101100011111010011111 ;
        654: q <= 32'b00111110000110010010100100100100 ;
        655: q <= 32'b10111110000010011001011010100100 ;
        656: q <= 32'b00111101000110010011100000110100 ;
        657: q <= 32'b10111100100111100001101110111100 ;
        658: q <= 32'b10111101000101100010101101110010 ;
        659: q <= 32'b00111101110100101101101010011001 ;
        660: q <= 32'b00111101100111100010011001110011 ;
        661: q <= 32'b00111100110110100101000101100000 ;
        662: q <= 32'b10111101110010011011001111011101 ;
        663: q <= 32'b10111110001011000100011000011100 ;
        664: q <= 32'b00111101110011101000001100001011 ;
        665: q <= 32'b00111101100000101111010000011100 ;
        666: q <= 32'b00111101001010110111011010010110 ;
        667: q <= 32'b10111101000100011110110111011000 ;
        668: q <= 32'b00111101000001100100100011111010 ;
        669: q <= 32'b10111101100101100101000010110010 ;
        670: q <= 32'b00111101101110011000000010110100 ;
        671: q <= 32'b10111101111001000011000100010000 ;
        672: q <= 32'b00111101110000011010100110100000 ;
        673: q <= 32'b00111101011111010111001010110000 ;
        674: q <= 32'b10111101101011010100101110011011 ;
        675: q <= 32'b00111011100100000001001101100011 ;
        676: q <= 32'b10111101110101001101001110010101 ;
        677: q <= 32'b10111101100110110000010110111101 ;
        678: q <= 32'b10111101110101011111100100111011 ;
        679: q <= 32'b10111101100111100100111110011110 ;
        680: q <= 32'b00111110000101000100000011100011 ;
        681: q <= 32'b00111101010011100100110010001010 ;
        682: q <= 32'b00111110000101011111010011101111 ;
        683: q <= 32'b10111101010011110010011111001110 ;
        684: q <= 32'b10111101100001010010101100011111 ;
        685: q <= 32'b10111101110111001010000100111101 ;
        686: q <= 32'b00111101101000110101000100101000 ;
        687: q <= 32'b00111101100011000011100000001000 ;
        688: q <= 32'b10111101111101010011111111011101 ;
        689: q <= 32'b10111101011111100000100011001110 ;
        690: q <= 32'b00111101000111101011011000000010 ;
        691: q <= 32'b00111100001110000010000010100101 ;
        692: q <= 32'b10111101000101000100010000000111 ;
        693: q <= 32'b00111101001001101001110111100011 ;
        694: q <= 32'b10111101000100010000111001011111 ;
        695: q <= 32'b00111100111100001111100010101110 ;
        696: q <= 32'b00111110000110101100000110011000 ;
        697: q <= 32'b10111101101111011110100001100110 ;
        698: q <= 32'b00111101101111110011100011010100 ;
        699: q <= 32'b00111101110101000111101111011101 ;
        700: q <= 32'b00111101100110011101011110011111 ;
        701: q <= 32'b10111010010001000111010010001111 ;
        702: q <= 32'b10111101010000110111001011101110 ;
        703: q <= 32'b10111101100111000100011000010110 ;
        704: q <= 32'b10111101010111110000010101100110 ;
        705: q <= 32'b10111101000101010000100100000010 ;
        706: q <= 32'b00111110001101101001101110000000 ;
        707: q <= 32'b10111100101001010011000100101101 ;
        708: q <= 32'b00111110000110101000110110101110 ;
        709: q <= 32'b10111100100110111111001100001000 ;
        710: q <= 32'b10111101110101001111111101111010 ;
        711: q <= 32'b00111010000000100100110100000100 ;
        712: q <= 32'b00111101001001000110011100110001 ;
        713: q <= 32'b10111101101100000001001011010001 ;
        714: q <= 32'b10111100100110101000101101100011 ;
        715: q <= 32'b00111101011011001101010100010010 ;
        716: q <= 32'b00111101011000011010110000010101 ;
        717: q <= 32'b10111100111011000011111101111110 ;
        718: q <= 32'b10111101011101101010110100011100 ;
        719: q <= 32'b10111100000110111100001100000000 ;
        720: q <= 32'b00111101100011011101100111110010 ;
        721: q <= 32'b00111110011000010011110111000000 ;
        722: q <= 32'b00111110000100001001101111000101 ;
        723: q <= 32'b10111101100001100111001111010111 ;
        724: q <= 32'b00111101111101110000010110110110 ;
        725: q <= 32'b00111110000100001100001110000100 ;
        726: q <= 32'b00111101101100010011110111100100 ;
        727: q <= 32'b00111100100010010000001000101000 ;
        728: q <= 32'b10111101000000011011101111001110 ;
        729: q <= 32'b00111101111110011001011010010010 ;
        730: q <= 32'b00111010110111100101011010000010 ;
        731: q <= 32'b00111101000101011010101010100110 ;
        732: q <= 32'b00111100111001011111101110001010 ;
        733: q <= 32'b10111101010101100011111100110010 ;
        734: q <= 32'b00111101110110111101000011110100 ;
        735: q <= 32'b10111101000101000001101100000010 ;
        736: q <= 32'b10111101011101100111001010011111 ;
        737: q <= 32'b00111101100010111100110001001100 ;
        738: q <= 32'b00111101010010110111101110101011 ;
        739: q <= 32'b00111101100001001110001110010101 ;
        740: q <= 32'b10111101011010110000100000011010 ;
        741: q <= 32'b00111110000011111110011000110101 ;
        742: q <= 32'b00111011011011111000010001010101 ;
        743: q <= 32'b00111100111100100010101101011101 ;
        744: q <= 32'b00000000000000000000000000000000 ;
        745: q <= 32'b00000000000000000000000000000000 ;
        746: q <= 32'b00000000000000000000000000000000 ;
        747: q <= 32'b00000000000000000000000000000000 ;
        748: q <= 32'b00000000000000000000000000000000 ;
        749: q <= 32'b00000000000000000000000000000000 ;
        750: q <= 32'b00000000000000000000000000000000 ;
        751: q <= 32'b00000000000000000000000000000000 ;
        752: q <= 32'b00000000000000000000000000000000 ;
        753: q <= 32'b00000000000000000000000000000000 ;
        754: q <= 32'b00000000000000000000000000000000 ;
        755: q <= 32'b00000000000000000000000000000000 ;
        756: q <= 32'b00000000000000000000000000000000 ;
        757: q <= 32'b00000000000000000000000000000000 ;
        758: q <= 32'b00000000000000000000000000000000 ;
        759: q <= 32'b00000000000000000000000000000000 ;
        760: q <= 32'b00000000000000000000000000000000 ;
        761: q <= 32'b00000000000000000000000000000000 ;
        762: q <= 32'b00000000000000000000000000000000 ;
        763: q <= 32'b00000000000000000000000000000000 ;
        764: q <= 32'b00000000000000000000000000000000 ;
        765: q <= 32'b00000000000000000000000000000000 ;
        766: q <= 32'b00000000000000000000000000000000 ;
        767: q <= 32'b00000000000000000000000000000000 ;
        768: q <= 32'b10111101111001101100000001110001 ;
        769: q <= 32'b00111101011000100001000001000010 ;
        770: q <= 32'b00111101100111101100111110111110 ;
        771: q <= 32'b00111101011010111001111011101001 ;
        772: q <= 32'b00111100100000001010000100110110 ;
        773: q <= 32'b00111100001000000001100010001001 ;
        774: q <= 32'b00111101001010110000101110110110 ;
        775: q <= 32'b00111101001001000101110111010010 ;
        776: q <= 32'b00111101011100010110001011111111 ;
        777: q <= 32'b00111101100110000001111101000000 ;
        778: q <= 32'b10111101000100010101111000101111 ;
        779: q <= 32'b10111101011110010111011110111001 ;
        780: q <= 32'b00111100110100000111001111110000 ;
        781: q <= 32'b10111101110000011000111001110000 ;
        782: q <= 32'b00111101000111110101001000000000 ;
        783: q <= 32'b10111101001110111000010101100001 ;
        784: q <= 32'b00111100101110011010000101111000 ;
        785: q <= 32'b00111101110001001100011011000101 ;
        786: q <= 32'b10111101100110101111000010011101 ;
        787: q <= 32'b00111101011010101111011001101110 ;
        788: q <= 32'b10111101100010011100010101001010 ;
        789: q <= 32'b10111101100011000101101100100110 ;
        790: q <= 32'b10111101010111101011110011011011 ;
        791: q <= 32'b10111101010010110000011010111001 ;
        792: q <= 32'b10111101101100011001010100011101 ;
        793: q <= 32'b10111100111001111001011010111001 ;
        794: q <= 32'b10111101011011001001001001111010 ;
        795: q <= 32'b10111100110101110010110010010001 ;
        796: q <= 32'b10111101111001111101000010000001 ;
        797: q <= 32'b00111101100010001100111000100111 ;
        798: q <= 32'b10111101110000001110100000011000 ;
        799: q <= 32'b00111101000001111010011011001001 ;
        800: q <= 32'b00111101010100111011001000010011 ;
        801: q <= 32'b10111100000100011110011111011100 ;
        802: q <= 32'b00111101101011110110101000101101 ;
        803: q <= 32'b10111101010000110011010011110011 ;
        804: q <= 32'b10111101001111111001111110001010 ;
        805: q <= 32'b10111101100111111010010100010011 ;
        806: q <= 32'b00111101001001110110000110100111 ;
        807: q <= 32'b00111101011000010010000001010110 ;
        808: q <= 32'b10111101000101111000001110010010 ;
        809: q <= 32'b10111101010011001100110000001100 ;
        810: q <= 32'b00111101100011110110000000100011 ;
        811: q <= 32'b00111101000110000101111100111101 ;
        812: q <= 32'b10111100101010011000000111111010 ;
        813: q <= 32'b10111100011010110011111100110110 ;
        814: q <= 32'b00111101101110100111001000011011 ;
        815: q <= 32'b10111101100011010100010100010110 ;
        816: q <= 32'b10111101100000110011100000111100 ;
        817: q <= 32'b10111101000011100000010010111110 ;
        818: q <= 32'b10111011011001111011010001000011 ;
        819: q <= 32'b00111101011100100001100111001110 ;
        820: q <= 32'b10111101000001111111110110100001 ;
        821: q <= 32'b10111101000001000011011010111011 ;
        822: q <= 32'b10111011100111101101101000100111 ;
        823: q <= 32'b00111101001010110100001110100111 ;
        824: q <= 32'b00111101100001011100011001100001 ;
        825: q <= 32'b10111101100010011100111010001010 ;
        826: q <= 32'b00111100110100110011110110100110 ;
        827: q <= 32'b00111100100111111000101000111011 ;
        828: q <= 32'b00111011000100000110101000000111 ;
        829: q <= 32'b00111100100000010111111000010110 ;
        830: q <= 32'b00111101100100011001100110001010 ;
        831: q <= 32'b00111011000011010010101100100101 ;
        832: q <= 32'b10111101101010011000111101000010 ;
        833: q <= 32'b10111101000000010110010111001110 ;
        834: q <= 32'b10111101000100101111100111111011 ;
        835: q <= 32'b10111101010000011000011100111011 ;
        836: q <= 32'b00111101101001000110010100101100 ;
        837: q <= 32'b10111100111101101111000001110011 ;
        838: q <= 32'b10111101100111110101010100101111 ;
        839: q <= 32'b10111101011010001111101000100111 ;
        840: q <= 32'b10111101100001110010111011100010 ;
        841: q <= 32'b00111101000110100100001011010101 ;
        842: q <= 32'b10111101010100010101110011110000 ;
        843: q <= 32'b00111100111010101111010001011001 ;
        844: q <= 32'b00111101001010010110100011000011 ;
        845: q <= 32'b00111100100011001110101011101100 ;
        846: q <= 32'b10111101101001010010101110000111 ;
        847: q <= 32'b10111100001011010110100001001101 ;
        848: q <= 32'b10111101100101101111010010011110 ;
        849: q <= 32'b10111100100010110101010011001100 ;
        850: q <= 32'b00111101100110111111110011111000 ;
        851: q <= 32'b10111101110001100000011110011011 ;
        852: q <= 32'b00111100111001111110011010010001 ;
        853: q <= 32'b10111101110101000111011010111000 ;
        854: q <= 32'b00111101101110010001100010011100 ;
        855: q <= 32'b00111101101100101101110101100111 ;
        856: q <= 32'b00111100011001100001011100101010 ;
        857: q <= 32'b10111010111011110110010110000100 ;
        858: q <= 32'b10111100101010111101100011111100 ;
        859: q <= 32'b10111101000100101010111001010010 ;
        860: q <= 32'b10111100100010100001001100100011 ;
        861: q <= 32'b00111101100111101111100100001010 ;
        862: q <= 32'b00111100101011001100110011001011 ;
        863: q <= 32'b10111101010010110111010101111010 ;
        864: q <= 32'b10111101001101110100101110111110 ;
        865: q <= 32'b10111101001001111110010001101111 ;
        866: q <= 32'b10111101101000000101111101011101 ;
        867: q <= 32'b10111010010110011011110001101110 ;
        868: q <= 32'b10111100000010110000001111100100 ;
        869: q <= 32'b10111100111100100000111010110110 ;
        870: q <= 32'b10111101100010100001001101100110 ;
        871: q <= 32'b00111100011001101011110100010101 ;
        872: q <= 32'b00000000000000000000000000000000 ;
        873: q <= 32'b00000000000000000000000000000000 ;
        874: q <= 32'b00000000000000000000000000000000 ;
        875: q <= 32'b00000000000000000000000000000000 ;
        876: q <= 32'b00000000000000000000000000000000 ;
        877: q <= 32'b00000000000000000000000000000000 ;
        878: q <= 32'b00000000000000000000000000000000 ;
        879: q <= 32'b00000000000000000000000000000000 ;
        880: q <= 32'b00000000000000000000000000000000 ;
        881: q <= 32'b00000000000000000000000000000000 ;
        882: q <= 32'b00000000000000000000000000000000 ;
        883: q <= 32'b00000000000000000000000000000000 ;
        884: q <= 32'b00000000000000000000000000000000 ;
        885: q <= 32'b00000000000000000000000000000000 ;
        886: q <= 32'b00000000000000000000000000000000 ;
        887: q <= 32'b00000000000000000000000000000000 ;
        888: q <= 32'b00000000000000000000000000000000 ;
        889: q <= 32'b00000000000000000000000000000000 ;
        890: q <= 32'b00000000000000000000000000000000 ;
        891: q <= 32'b00000000000000000000000000000000 ;
        892: q <= 32'b00000000000000000000000000000000 ;
        893: q <= 32'b00000000000000000000000000000000 ;
        894: q <= 32'b00000000000000000000000000000000 ;
        895: q <= 32'b00000000000000000000000000000000 ;
        896: q <= 32'b10111010100001110110111100111001 ;
        897: q <= 32'b10111101110011001101111110011110 ;
        898: q <= 32'b00111100001111010011010110100010 ;
        899: q <= 32'b10111101111011010010001010001001 ;
        900: q <= 32'b10111011110110000101110100001011 ;
        901: q <= 32'b00111101100000010111111101110100 ;
        902: q <= 32'b00111101000110101100011110110100 ;
        903: q <= 32'b10111101100001110000010100011001 ;
        904: q <= 32'b00111101001000101011100101010011 ;
        905: q <= 32'b10111100100010110001000000011111 ;
        906: q <= 32'b10111100110001100000100010111011 ;
        907: q <= 32'b10111101100001101111011001000100 ;
        908: q <= 32'b00111101101111001010101111001101 ;
        909: q <= 32'b10111101110011000011011111101001 ;
        910: q <= 32'b10111101000100111110101011101011 ;
        911: q <= 32'b10111101101101000100001000001101 ;
        912: q <= 32'b10111101011010001000001000101000 ;
        913: q <= 32'b10111100111001110100001001101100 ;
        914: q <= 32'b00111101001111110111110001000001 ;
        915: q <= 32'b10111101001110000101111010000101 ;
        916: q <= 32'b10111101100001000011011110110011 ;
        917: q <= 32'b10111101110000011111010001000101 ;
        918: q <= 32'b10111100101100100111110111101110 ;
        919: q <= 32'b10111101101101011110100001100110 ;
        920: q <= 32'b00111101100101100010010101011001 ;
        921: q <= 32'b10111010111100010010110001010010 ;
        922: q <= 32'b10111110000000100001110111100110 ;
        923: q <= 32'b10111101101011001100110010011010 ;
        924: q <= 32'b10111101100100000110111110001110 ;
        925: q <= 32'b10111101110101010010000111111100 ;
        926: q <= 32'b00111101011011010111111000010100 ;
        927: q <= 32'b10111100100101101100010100000000 ;
        928: q <= 32'b00111101011010011000100001111001 ;
        929: q <= 32'b10111101100101100110101001001111 ;
        930: q <= 32'b10111101101110001011001110111000 ;
        931: q <= 32'b00111101011010101000000101010110 ;
        932: q <= 32'b00111101010111101010111011011101 ;
        933: q <= 32'b00111011110101110001001010100000 ;
        934: q <= 32'b10111100000010001101110101110110 ;
        935: q <= 32'b10111100001010110111000010110111 ;
        936: q <= 32'b10111100100111010011000000110100 ;
        937: q <= 32'b10111101001001011100100011101001 ;
        938: q <= 32'b00111100110110010000111111100011 ;
        939: q <= 32'b10111101000101011110110011101111 ;
        940: q <= 32'b10111100110011010011000100001001 ;
        941: q <= 32'b00111101101111111010110111100111 ;
        942: q <= 32'b00111101101101010011100000010100 ;
        943: q <= 32'b00111101100011011010100111111111 ;
        944: q <= 32'b10111100000111101011011101100101 ;
        945: q <= 32'b00111101101110101001011000000101 ;
        946: q <= 32'b00111101011100010100001110000110 ;
        947: q <= 32'b10111100000001110101111100100000 ;
        948: q <= 32'b10111011110110111101011111000100 ;
        949: q <= 32'b00111101000001100101000111000100 ;
        950: q <= 32'b10111101111000000101001110101111 ;
        951: q <= 32'b10111101100000110100101000011101 ;
        952: q <= 32'b00111101001110101011001101110110 ;
        953: q <= 32'b10111101100011010110001111001101 ;
        954: q <= 32'b00111101000010011111100000111101 ;
        955: q <= 32'b00111100000101100101111110110100 ;
        956: q <= 32'b10111101011101100101001000001000 ;
        957: q <= 32'b10111100101110101010111010101001 ;
        958: q <= 32'b00111101000100011100101000101101 ;
        959: q <= 32'b10111101011101001011110010011101 ;
        960: q <= 32'b00111101011001110110111110111011 ;
        961: q <= 32'b00111101110111101001110111011111 ;
        962: q <= 32'b00111101011100100000110100001010 ;
        963: q <= 32'b10111101110010111000010100110010 ;
        964: q <= 32'b10111101100000101010001101001111 ;
        965: q <= 32'b10111100011111111100000001000001 ;
        966: q <= 32'b10111010111010110001100010101001 ;
        967: q <= 32'b00111100111000110000101011100010 ;
        968: q <= 32'b00111101001111011000110101000101 ;
        969: q <= 32'b10111101011111111101100011111110 ;
        970: q <= 32'b00111100010011001000000111101110 ;
        971: q <= 32'b10111101100000000000001111000010 ;
        972: q <= 32'b10111101101001001110110011010001 ;
        973: q <= 32'b00111100100011101111011010000110 ;
        974: q <= 32'b10111101111001000000001110011100 ;
        975: q <= 32'b10111010101010010110111110100110 ;
        976: q <= 32'b00111100101011001001110101010110 ;
        977: q <= 32'b00111101100100101101111101100110 ;
        978: q <= 32'b00111100010110011111010010001001 ;
        979: q <= 32'b10111101110100100110101011010110 ;
        980: q <= 32'b00111100111110110010100000111011 ;
        981: q <= 32'b00111101001110100011110110110111 ;
        982: q <= 32'b00111101110000101100001101100011 ;
        983: q <= 32'b10111101101000100001000001000111 ;
        984: q <= 32'b10111101101111111100111101001011 ;
        985: q <= 32'b10111011111010101000111000101111 ;
        986: q <= 32'b00111101101111110110101001111101 ;
        987: q <= 32'b00111101000101100011111011101110 ;
        988: q <= 32'b00111100001001011000000010011011 ;
        989: q <= 32'b10111101011100100011011101001010 ;
        990: q <= 32'b10111100101110001101000011000100 ;
        991: q <= 32'b10111101010001010100001110001011 ;
        992: q <= 32'b00111101100000110011010111111011 ;
        993: q <= 32'b10111100100010010101100111001010 ;
        994: q <= 32'b10111101000001101011100011111011 ;
        995: q <= 32'b00111101010110101111100101010101 ;
        996: q <= 32'b10111100010001010000111001110011 ;
        997: q <= 32'b00111101110000001100000000011100 ;
        998: q <= 32'b10111101001110110110010010111100 ;
        999: q <= 32'b10111100101000111111010100011011 ;
        1000: q <= 32'b00000000000000000000000000000000 ;
        1001: q <= 32'b00000000000000000000000000000000 ;
        1002: q <= 32'b00000000000000000000000000000000 ;
        1003: q <= 32'b00000000000000000000000000000000 ;
        1004: q <= 32'b00000000000000000000000000000000 ;
        1005: q <= 32'b00000000000000000000000000000000 ;
        1006: q <= 32'b00000000000000000000000000000000 ;
        1007: q <= 32'b00000000000000000000000000000000 ;
        1008: q <= 32'b00000000000000000000000000000000 ;
        1009: q <= 32'b00000000000000000000000000000000 ;
        1010: q <= 32'b00000000000000000000000000000000 ;
        1011: q <= 32'b00000000000000000000000000000000 ;
        1012: q <= 32'b00000000000000000000000000000000 ;
        1013: q <= 32'b00000000000000000000000000000000 ;
        1014: q <= 32'b00000000000000000000000000000000 ;
        1015: q <= 32'b00000000000000000000000000000000 ;
        1016: q <= 32'b00000000000000000000000000000000 ;
        1017: q <= 32'b00000000000000000000000000000000 ;
        1018: q <= 32'b00000000000000000000000000000000 ;
        1019: q <= 32'b00000000000000000000000000000000 ;
        1020: q <= 32'b00000000000000000000000000000000 ;
        1021: q <= 32'b00000000000000000000000000000000 ;
        1022: q <= 32'b00000000000000000000000000000000 ;
        1023: q <= 32'b00000000000000000000000000000000 ;
        1024: q <= 32'b00111100100111010100100011110001 ;
        1025: q <= 32'b10111101000010101001101001011111 ;
        1026: q <= 32'b10111100111000011101000011101100 ;
        1027: q <= 32'b10111110000001100101000110011101 ;
        1028: q <= 32'b00111100000111001111110000111000 ;
        1029: q <= 32'b10111101101010010110100111000001 ;
        1030: q <= 32'b10111101100011001111111011000010 ;
        1031: q <= 32'b10111101001110110010000001101111 ;
        1032: q <= 32'b10111100111100000111000101010010 ;
        1033: q <= 32'b00111110000000010100110111010110 ;
        1034: q <= 32'b10111110000000101111001000101000 ;
        1035: q <= 32'b00111101010010001111010110011011 ;
        1036: q <= 32'b00111101111000000010100110000110 ;
        1037: q <= 32'b00111100101001001000000111100110 ;
        1038: q <= 32'b00111101110110110110011110100010 ;
        1039: q <= 32'b10111101100110101010100010001001 ;
        1040: q <= 32'b10111100111101010111101101111000 ;
        1041: q <= 32'b00111101101011010110000001001101 ;
        1042: q <= 32'b10111101111110110101111100101011 ;
        1043: q <= 32'b10111011111011000100001000111011 ;
        1044: q <= 32'b10111100111000000000111111101011 ;
        1045: q <= 32'b10111101101100100111011100000110 ;
        1046: q <= 32'b00111101010100100110111100111111 ;
        1047: q <= 32'b00111100101010100110001111110000 ;
        1048: q <= 32'b00111101100011000110111110100111 ;
        1049: q <= 32'b00111100101111110010111100101000 ;
        1050: q <= 32'b10111101010101000011000101011110 ;
        1051: q <= 32'b10111100010011010001011110101001 ;
        1052: q <= 32'b00111110000100111101000011001101 ;
        1053: q <= 32'b10111110000111100100111000101111 ;
        1054: q <= 32'b10111101111100011111001101010010 ;
        1055: q <= 32'b10111101010000100001111011100111 ;
        1056: q <= 32'b00111100000101100011111101001101 ;
        1057: q <= 32'b00111100010100101101010001111000 ;
        1058: q <= 32'b00111101011001000101100011110101 ;
        1059: q <= 32'b00111110000000000010111001010100 ;
        1060: q <= 32'b10111101111110011001111001010111 ;
        1061: q <= 32'b10111011110110011100111100011000 ;
        1062: q <= 32'b10111011100110011001001110010011 ;
        1063: q <= 32'b00111011110100010010100010110111 ;
        1064: q <= 32'b10111101100110110001110010001100 ;
        1065: q <= 32'b00111101110011100110111101101110 ;
        1066: q <= 32'b00111101100110100100010001111000 ;
        1067: q <= 32'b00111100111111011111011001010010 ;
        1068: q <= 32'b10111101010000101001111110011111 ;
        1069: q <= 32'b00111101010001010000001011110101 ;
        1070: q <= 32'b10111101101101111010001101100000 ;
        1071: q <= 32'b10111100101100011101110100100011 ;
        1072: q <= 32'b10111101111001100101100011011100 ;
        1073: q <= 32'b10111101101010110110011010110000 ;
        1074: q <= 32'b00111101010000101001000001110000 ;
        1075: q <= 32'b10111011111010100010100001100110 ;
        1076: q <= 32'b10111101111101011010110000111001 ;
        1077: q <= 32'b10111100100001110101000111111000 ;
        1078: q <= 32'b00111101100110000100011101100010 ;
        1079: q <= 32'b10111101110010001101001110101100 ;
        1080: q <= 32'b00111101101000100111001010011011 ;
        1081: q <= 32'b00111100001110111011111000101111 ;
        1082: q <= 32'b10111011111000001010010111110001 ;
        1083: q <= 32'b10111101011110111110111111011011 ;
        1084: q <= 32'b10111101000010110101101111011010 ;
        1085: q <= 32'b10111101100001010111010111101000 ;
        1086: q <= 32'b00111011100110001110111100000100 ;
        1087: q <= 32'b00111110000000000110101100101011 ;
        1088: q <= 32'b00111101110100000011011111010111 ;
        1089: q <= 32'b10111011100001110000110101011000 ;
        1090: q <= 32'b10111100101110000011000100011101 ;
        1091: q <= 32'b00111101101111101111000001110010 ;
        1092: q <= 32'b00111110000010100101100000100000 ;
        1093: q <= 32'b00111100100001111011110110001100 ;
        1094: q <= 32'b10111101011101010011110111110101 ;
        1095: q <= 32'b10111101111111010100011101001100 ;
        1096: q <= 32'b10111101010101011011101000101110 ;
        1097: q <= 32'b00111110000001111011110110100010 ;
        1098: q <= 32'b10111101101100110010010010101111 ;
        1099: q <= 32'b00111101101110110011100000011101 ;
        1100: q <= 32'b10111101001011101111010110101111 ;
        1101: q <= 32'b00111100111001100000001110010001 ;
        1102: q <= 32'b10111100111001000010010100110111 ;
        1103: q <= 32'b10111100101011011101100001001111 ;
        1104: q <= 32'b10111100010001111000111101100101 ;
        1105: q <= 32'b00111101110000001110111000100010 ;
        1106: q <= 32'b10111100100011001010010100011000 ;
        1107: q <= 32'b10111110000110101001000100000010 ;
        1108: q <= 32'b00111011011001110010010100011001 ;
        1109: q <= 32'b10111101101000111001001100111110 ;
        1110: q <= 32'b10111100010000001000110011011011 ;
        1111: q <= 32'b00111101001110110110001001001011 ;
        1112: q <= 32'b00111011101101111000101011101100 ;
        1113: q <= 32'b10111101011101011101010100000111 ;
        1114: q <= 32'b10111100111100001101101000101001 ;
        1115: q <= 32'b10111101111101111101000010101001 ;
        1116: q <= 32'b00111101101001010000111000001101 ;
        1117: q <= 32'b00111101001100100000111110110111 ;
        1118: q <= 32'b00111110000010000101100001001011 ;
        1119: q <= 32'b00111100000111110110000111101111 ;
        1120: q <= 32'b10111101100000110111000110010011 ;
        1121: q <= 32'b00111100111000111100010111110001 ;
        1122: q <= 32'b10111101110100100110011001101111 ;
        1123: q <= 32'b10111101010110001001010101011101 ;
        1124: q <= 32'b10111101001001101000010011000010 ;
        1125: q <= 32'b10111100100111010000000000110101 ;
        1126: q <= 32'b00111101101110011001110100110111 ;
        1127: q <= 32'b00111101001001000101111010011111 ;
        1128: q <= 32'b00000000000000000000000000000000 ;
        1129: q <= 32'b00000000000000000000000000000000 ;
        1130: q <= 32'b00000000000000000000000000000000 ;
        1131: q <= 32'b00000000000000000000000000000000 ;
        1132: q <= 32'b00000000000000000000000000000000 ;
        1133: q <= 32'b00000000000000000000000000000000 ;
        1134: q <= 32'b00000000000000000000000000000000 ;
        1135: q <= 32'b00000000000000000000000000000000 ;
        1136: q <= 32'b00000000000000000000000000000000 ;
        1137: q <= 32'b00000000000000000000000000000000 ;
        1138: q <= 32'b00000000000000000000000000000000 ;
        1139: q <= 32'b00000000000000000000000000000000 ;
        1140: q <= 32'b00000000000000000000000000000000 ;
        1141: q <= 32'b00000000000000000000000000000000 ;
        1142: q <= 32'b00000000000000000000000000000000 ;
        1143: q <= 32'b00000000000000000000000000000000 ;
        1144: q <= 32'b00000000000000000000000000000000 ;
        1145: q <= 32'b00000000000000000000000000000000 ;
        1146: q <= 32'b00000000000000000000000000000000 ;
        1147: q <= 32'b00000000000000000000000000000000 ;
        1148: q <= 32'b00000000000000000000000000000000 ;
        1149: q <= 32'b00000000000000000000000000000000 ;
        1150: q <= 32'b00000000000000000000000000000000 ;
        1151: q <= 32'b00000000000000000000000000000000 ;
        1152: q <= 32'b00111110000000010011110100011101 ;
        1153: q <= 32'b10111101100010001101110110000010 ;
        1154: q <= 32'b10111101110001101011011000000010 ;
        1155: q <= 32'b10111011110110101110010101001100 ;
        1156: q <= 32'b00111101100111000110000101100111 ;
        1157: q <= 32'b00111101000010011110100010001110 ;
        1158: q <= 32'b00111101110000000000010011101000 ;
        1159: q <= 32'b10111110001011001001100011101100 ;
        1160: q <= 32'b00111110001011011011011011111001 ;
        1161: q <= 32'b10111101101010100110100000100110 ;
        1162: q <= 32'b10111101101001101100110100101110 ;
        1163: q <= 32'b10111101110111000101100100100100 ;
        1164: q <= 32'b00111101101111011111111000011100 ;
        1165: q <= 32'b10111101111001001110000101001110 ;
        1166: q <= 32'b10111101111100011110100010010100 ;
        1167: q <= 32'b00111101100010110010001001001111 ;
        1168: q <= 32'b00111101101011111101011001110111 ;
        1169: q <= 32'b10111101010101001100110001111001 ;
        1170: q <= 32'b00111100001010011010001111000100 ;
        1171: q <= 32'b00111101000001010101010101110111 ;
        1172: q <= 32'b00111101111111011010000010010000 ;
        1173: q <= 32'b00111011110101100011010010001100 ;
        1174: q <= 32'b10111100111111100110010110011110 ;
        1175: q <= 32'b10111101011101011100001001110010 ;
        1176: q <= 32'b10111100101011000101100001010111 ;
        1177: q <= 32'b00111010110100011000110101101010 ;
        1178: q <= 32'b10111101100100011010101011001000 ;
        1179: q <= 32'b00111100110101111111011010001100 ;
        1180: q <= 32'b10111100000101001000111011000111 ;
        1181: q <= 32'b00111101010110000111110010111111 ;
        1182: q <= 32'b10111101011101100001110010100110 ;
        1183: q <= 32'b10111100011111101010011101011010 ;
        1184: q <= 32'b10111100110011110100100001010100 ;
        1185: q <= 32'b10111101100101000000110010101010 ;
        1186: q <= 32'b10111100011111010001000000001001 ;
        1187: q <= 32'b10111100011111100010000011001000 ;
        1188: q <= 32'b00111101100111000100101011000000 ;
        1189: q <= 32'b00111100110010100100001001011101 ;
        1190: q <= 32'b10111101110001111110111110100111 ;
        1191: q <= 32'b10111101100001111011001110000100 ;
        1192: q <= 32'b00111110000001011010110100100110 ;
        1193: q <= 32'b00111101101010011000000100011110 ;
        1194: q <= 32'b10111010100001011110010111000110 ;
        1195: q <= 32'b10111101111001001110000111100000 ;
        1196: q <= 32'b00111100001010001010001001110001 ;
        1197: q <= 32'b10111101111110100101110010101100 ;
        1198: q <= 32'b10111101000101100101111111111111 ;
        1199: q <= 32'b00111101001001011011101100001011 ;
        1200: q <= 32'b00111101001111101101100000100111 ;
        1201: q <= 32'b00111110000001101001100101010010 ;
        1202: q <= 32'b00111100000101111000000101111011 ;
        1203: q <= 32'b10111101001110001000000000011001 ;
        1204: q <= 32'b10111101111010110100010011101010 ;
        1205: q <= 32'b00111100101000101111111110110101 ;
        1206: q <= 32'b00111100110110010010010110110100 ;
        1207: q <= 32'b00111100100100100011010100111001 ;
        1208: q <= 32'b00111101100010110111011010110010 ;
        1209: q <= 32'b00111101011110101001000000100011 ;
        1210: q <= 32'b00111101110111101000110010100000 ;
        1211: q <= 32'b00111101000011110111111010100111 ;
        1212: q <= 32'b00111101101100010111010001001000 ;
        1213: q <= 32'b10111101101110011111001000111011 ;
        1214: q <= 32'b00111011110000011100110000100100 ;
        1215: q <= 32'b00111101000110111101011101110010 ;
        1216: q <= 32'b00111100000100000101010001001100 ;
        1217: q <= 32'b10111110000001011101101000000110 ;
        1218: q <= 32'b00111101011000101000111010010000 ;
        1219: q <= 32'b10111100111010111011111001111111 ;
        1220: q <= 32'b00111100100100001011110010101100 ;
        1221: q <= 32'b00111101011011110111010010000110 ;
        1222: q <= 32'b10111100111110001111011100101001 ;
        1223: q <= 32'b10111101100101101100000100100101 ;
        1224: q <= 32'b10111101010011010100110110011011 ;
        1225: q <= 32'b10111110000110100101100111100100 ;
        1226: q <= 32'b10111001101110011100101101101001 ;
        1227: q <= 32'b00111101100110001000000000000010 ;
        1228: q <= 32'b00111011111111010011110111000010 ;
        1229: q <= 32'b00111101101111100110111010001000 ;
        1230: q <= 32'b00111100111100011010111001100100 ;
        1231: q <= 32'b00111101100011100110000001000001 ;
        1232: q <= 32'b10111101000010001011001000010111 ;
        1233: q <= 32'b10111011100111001100100100010101 ;
        1234: q <= 32'b10111101011011110110000010101010 ;
        1235: q <= 32'b00111101011110000110101100100010 ;
        1236: q <= 32'b10111101011101110000110010011101 ;
        1237: q <= 32'b10111101001110100101010110001101 ;
        1238: q <= 32'b10111101011000000100101100011100 ;
        1239: q <= 32'b00111101010001010011110100010110 ;
        1240: q <= 32'b10111100100001010000111000101101 ;
        1241: q <= 32'b10111101011110001100111010100111 ;
        1242: q <= 32'b00111101001100000000011010100111 ;
        1243: q <= 32'b10111101011111111001000101111001 ;
        1244: q <= 32'b00111101010100001000111001100110 ;
        1245: q <= 32'b10111101011010111111011100001110 ;
        1246: q <= 32'b00111100110011001101101100101001 ;
        1247: q <= 32'b10111101100000010001110001011000 ;
        1248: q <= 32'b00111101111000001011110010101110 ;
        1249: q <= 32'b00111010111101000111001001101101 ;
        1250: q <= 32'b00111101101101011111110100101110 ;
        1251: q <= 32'b10111011000111010000110111001010 ;
        1252: q <= 32'b00111101011011101101001110011011 ;
        1253: q <= 32'b00111101010111010010110000011001 ;
        1254: q <= 32'b00111101100011111101001000101101 ;
        1255: q <= 32'b00111100110000010010111101101001 ;
        1256: q <= 32'b00000000000000000000000000000000 ;
        1257: q <= 32'b00000000000000000000000000000000 ;
        1258: q <= 32'b00000000000000000000000000000000 ;
        1259: q <= 32'b00000000000000000000000000000000 ;
        1260: q <= 32'b00000000000000000000000000000000 ;
        1261: q <= 32'b00000000000000000000000000000000 ;
        1262: q <= 32'b00000000000000000000000000000000 ;
        1263: q <= 32'b00000000000000000000000000000000 ;
        1264: q <= 32'b00000000000000000000000000000000 ;
        1265: q <= 32'b00000000000000000000000000000000 ;
        1266: q <= 32'b00000000000000000000000000000000 ;
        1267: q <= 32'b00000000000000000000000000000000 ;
        1268: q <= 32'b00000000000000000000000000000000 ;
        1269: q <= 32'b00000000000000000000000000000000 ;
        1270: q <= 32'b00000000000000000000000000000000 ;
        1271: q <= 32'b00000000000000000000000000000000 ;
        1272: q <= 32'b00000000000000000000000000000000 ;
        1273: q <= 32'b00000000000000000000000000000000 ;
        1274: q <= 32'b00000000000000000000000000000000 ;
        1275: q <= 32'b00000000000000000000000000000000 ;
        1276: q <= 32'b00000000000000000000000000000000 ;
        1277: q <= 32'b00000000000000000000000000000000 ;
        1278: q <= 32'b00000000000000000000000000000000 ;
        1279: q <= 32'b00000000000000000000000000000000 ;
        1280: q <= 32'b10111101000100111011100000101001 ;
        1281: q <= 32'b00111011000100111111100000000100 ;
        1282: q <= 32'b10111101110101000001100000010000 ;
        1283: q <= 32'b10111100001000011111110111110011 ;
        1284: q <= 32'b00111110000110111100111011001110 ;
        1285: q <= 32'b00111100100110100100111101110011 ;
        1286: q <= 32'b10111110010010101111101111011000 ;
        1287: q <= 32'b10111100100101110000100111011101 ;
        1288: q <= 32'b00111011101011011010000100011001 ;
        1289: q <= 32'b00111100011110111010101000111100 ;
        1290: q <= 32'b00111101111100110011011001000100 ;
        1291: q <= 32'b10111100111001111100100010100110 ;
        1292: q <= 32'b10111011110000011111011110001100 ;
        1293: q <= 32'b00111100000110001010011100100010 ;
        1294: q <= 32'b10111101100110110111101110000001 ;
        1295: q <= 32'b00111110000011101101100110110110 ;
        1296: q <= 32'b00111101011110010100010100110110 ;
        1297: q <= 32'b10111101100100011011110110001011 ;
        1298: q <= 32'b00111101000000001110110001001000 ;
        1299: q <= 32'b00111110000101000110010001010011 ;
        1300: q <= 32'b10111101101000100001100101010100 ;
        1301: q <= 32'b00111100000111000011111001100000 ;
        1302: q <= 32'b00111101100101001010010000101111 ;
        1303: q <= 32'b10111101101011111011001111111010 ;
        1304: q <= 32'b10111110001110000010101100000101 ;
        1305: q <= 32'b00111100100010000111101010101000 ;
        1306: q <= 32'b00111101010001101100111111111101 ;
        1307: q <= 32'b10111100111000110110001011010000 ;
        1308: q <= 32'b10111101111110010110001100000110 ;
        1309: q <= 32'b00111101110100001000010101110010 ;
        1310: q <= 32'b00111110000110111010001000111101 ;
        1311: q <= 32'b10111010101111101010011010110001 ;
        1312: q <= 32'b10111101010001111110110010111011 ;
        1313: q <= 32'b00111100010001110010101100110011 ;
        1314: q <= 32'b10111011110111000001101001000000 ;
        1315: q <= 32'b00111101101010101100111110000011 ;
        1316: q <= 32'b10111101010110011101110011101110 ;
        1317: q <= 32'b10111101100011001010011101110101 ;
        1318: q <= 32'b00111011001100100001100110110101 ;
        1319: q <= 32'b00111101000000111011110010101110 ;
        1320: q <= 32'b10111101101000110100000011100100 ;
        1321: q <= 32'b10111101001101111011010111110010 ;
        1322: q <= 32'b10111101000010110010011101010000 ;
        1323: q <= 32'b00111010010010111100001001100101 ;
        1324: q <= 32'b00111101111001011101001011001111 ;
        1325: q <= 32'b00111101111101011100101011001100 ;
        1326: q <= 32'b10111010011101100100100000111010 ;
        1327: q <= 32'b10111101111010100100110011000010 ;
        1328: q <= 32'b00111101101101110010000010011001 ;
        1329: q <= 32'b00111101100111000110010100101000 ;
        1330: q <= 32'b10111101101110011100101110110110 ;
        1331: q <= 32'b00111101101001101010011110001000 ;
        1332: q <= 32'b10111101100010111011010110001111 ;
        1333: q <= 32'b00111101000110100000111110001101 ;
        1334: q <= 32'b10111100100110001010100101100000 ;
        1335: q <= 32'b10111101100110000111101000100011 ;
        1336: q <= 32'b00111101010000110011001111010110 ;
        1337: q <= 32'b10111101100110010001000110101011 ;
        1338: q <= 32'b10111101101101000000101000100011 ;
        1339: q <= 32'b00111100110100110001100001001001 ;
        1340: q <= 32'b00111101011000000111110101110000 ;
        1341: q <= 32'b00111101000010001101000100111010 ;
        1342: q <= 32'b10111100111101011111011110111011 ;
        1343: q <= 32'b00111100000000101010010100110100 ;
        1344: q <= 32'b00111100001001111010001101010011 ;
        1345: q <= 32'b10111101101011100101000110101011 ;
        1346: q <= 32'b10111101010110011101011111111100 ;
        1347: q <= 32'b10111100111101011111000101110000 ;
        1348: q <= 32'b10111101010010111001001111110111 ;
        1349: q <= 32'b00111101011011011010011101110101 ;
        1350: q <= 32'b00111011000111011100110000111010 ;
        1351: q <= 32'b00111100000111000000000100100111 ;
        1352: q <= 32'b10111100001001100001101000000001 ;
        1353: q <= 32'b10111101110111110110010000010010 ;
        1354: q <= 32'b00111101100100000111110000001000 ;
        1355: q <= 32'b10111101001001000111010101100110 ;
        1356: q <= 32'b10111100100010110011100001001011 ;
        1357: q <= 32'b00111101010101111111111110111001 ;
        1358: q <= 32'b00111101100011011110011001101000 ;
        1359: q <= 32'b00111110001101111100111000100010 ;
        1360: q <= 32'b10111101111011111001110010111010 ;
        1361: q <= 32'b10111110000011001111100100011101 ;
        1362: q <= 32'b00111100111111011100011100010101 ;
        1363: q <= 32'b10111100000010100111011001110001 ;
        1364: q <= 32'b10111101011101011000000111110010 ;
        1365: q <= 32'b10111101010100100110100110010000 ;
        1366: q <= 32'b10111100101101011101110010110000 ;
        1367: q <= 32'b10111100000001100011101010010000 ;
        1368: q <= 32'b00111101011100011101000100110111 ;
        1369: q <= 32'b00111101000011010000010110011001 ;
        1370: q <= 32'b10111100111001110011010010100011 ;
        1371: q <= 32'b10111101000110000000100001111001 ;
        1372: q <= 32'b00111010111001111101010001011111 ;
        1373: q <= 32'b10111110000000111000111100001011 ;
        1374: q <= 32'b10111101100110010011110011011010 ;
        1375: q <= 32'b10111101000000001000000010010011 ;
        1376: q <= 32'b10111100100111100110110000000100 ;
        1377: q <= 32'b10111101110010000001001111000111 ;
        1378: q <= 32'b10111101101011100110000101010001 ;
        1379: q <= 32'b10111101101110100010011001001111 ;
        1380: q <= 32'b00111101011001111011011111011100 ;
        1381: q <= 32'b10111101100110101110101111110110 ;
        1382: q <= 32'b00111101100110010101100001110010 ;
        1383: q <= 32'b00111101011001011111101110010101 ;
        1384: q <= 32'b00000000000000000000000000000000 ;
        1385: q <= 32'b00000000000000000000000000000000 ;
        1386: q <= 32'b00000000000000000000000000000000 ;
        1387: q <= 32'b00000000000000000000000000000000 ;
        1388: q <= 32'b00000000000000000000000000000000 ;
        1389: q <= 32'b00000000000000000000000000000000 ;
        1390: q <= 32'b00000000000000000000000000000000 ;
        1391: q <= 32'b00000000000000000000000000000000 ;
        1392: q <= 32'b00000000000000000000000000000000 ;
        1393: q <= 32'b00000000000000000000000000000000 ;
        1394: q <= 32'b00000000000000000000000000000000 ;
        1395: q <= 32'b00000000000000000000000000000000 ;
        1396: q <= 32'b00000000000000000000000000000000 ;
        1397: q <= 32'b00000000000000000000000000000000 ;
        1398: q <= 32'b00000000000000000000000000000000 ;
        1399: q <= 32'b00000000000000000000000000000000 ;
        1400: q <= 32'b00000000000000000000000000000000 ;
        1401: q <= 32'b00000000000000000000000000000000 ;
        1402: q <= 32'b00000000000000000000000000000000 ;
        1403: q <= 32'b00000000000000000000000000000000 ;
        1404: q <= 32'b00000000000000000000000000000000 ;
        1405: q <= 32'b00000000000000000000000000000000 ;
        1406: q <= 32'b00000000000000000000000000000000 ;
        1407: q <= 32'b00000000000000000000000000000000 ;
        1408: q <= 32'b10111110000011101101100100011110 ;
        1409: q <= 32'b00111101001100111101100001000100 ;
        1410: q <= 32'b10111100000011101110000100001001 ;
        1411: q <= 32'b10111100000101111100001000000100 ;
        1412: q <= 32'b10111101110110110000000011001000 ;
        1413: q <= 32'b00111011101101111001111011101100 ;
        1414: q <= 32'b10111001100011100111100101111011 ;
        1415: q <= 32'b00111101100101011001101010000100 ;
        1416: q <= 32'b10111101000010000111101000100100 ;
        1417: q <= 32'b00111100000100010110110010100011 ;
        1418: q <= 32'b00111100010111110111011101100111 ;
        1419: q <= 32'b00111101101101000000100100011001 ;
        1420: q <= 32'b00111101001111111100100101110010 ;
        1421: q <= 32'b00111110000110100101011111110011 ;
        1422: q <= 32'b10111011101101001010110110011010 ;
        1423: q <= 32'b00111100110110001111101100111001 ;
        1424: q <= 32'b10111101000010000101110011010010 ;
        1425: q <= 32'b10111101001111010011111011100110 ;
        1426: q <= 32'b00111101001000000001110011000011 ;
        1427: q <= 32'b00111101000000111100101100000111 ;
        1428: q <= 32'b00111100101111110110001111010100 ;
        1429: q <= 32'b10111101110001001111100000000011 ;
        1430: q <= 32'b00111101110010101110011001001101 ;
        1431: q <= 32'b10111100101100111101111010100011 ;
        1432: q <= 32'b00111101011000011010000000001011 ;
        1433: q <= 32'b10111100111000111101011111010011 ;
        1434: q <= 32'b10111101111001111101111010111011 ;
        1435: q <= 32'b00111100101011101011000000111110 ;
        1436: q <= 32'b00111101110111000011100010011100 ;
        1437: q <= 32'b10111101100000110101111111001100 ;
        1438: q <= 32'b10111101101001010001000011011011 ;
        1439: q <= 32'b00111100101001001000100101001000 ;
        1440: q <= 32'b00111101100011000110111011100110 ;
        1441: q <= 32'b10111101100001001111000111000100 ;
        1442: q <= 32'b10111101010100100101010101000010 ;
        1443: q <= 32'b00111101011001000100000011000101 ;
        1444: q <= 32'b10111101010100101110110001111010 ;
        1445: q <= 32'b10111101000010101101000000110001 ;
        1446: q <= 32'b10111000101011111011100101011110 ;
        1447: q <= 32'b00111110000101001011100111011001 ;
        1448: q <= 32'b00111101110011010011000011001100 ;
        1449: q <= 32'b00111101001111101110000100111010 ;
        1450: q <= 32'b10111110001001110110100000001010 ;
        1451: q <= 32'b10111100000111010011010000100110 ;
        1452: q <= 32'b10111011101001111001011010110010 ;
        1453: q <= 32'b10111101000001110011000001011110 ;
        1454: q <= 32'b00111101001000001011011010010011 ;
        1455: q <= 32'b00111101011000001001111100101111 ;
        1456: q <= 32'b10111101100010001010010011001010 ;
        1457: q <= 32'b00111101011111011000011001101101 ;
        1458: q <= 32'b10111101010101000000001110001111 ;
        1459: q <= 32'b00111100110101101010101001010110 ;
        1460: q <= 32'b10111101100001111100010100000101 ;
        1461: q <= 32'b00111101101010101010101011111111 ;
        1462: q <= 32'b10111100111010101110010001110010 ;
        1463: q <= 32'b00111010101110011000001010101101 ;
        1464: q <= 32'b00111011111010010100100010010011 ;
        1465: q <= 32'b10111101101001010110000100110000 ;
        1466: q <= 32'b10111011110101010001111101101000 ;
        1467: q <= 32'b10111100100001110001000101001010 ;
        1468: q <= 32'b10111101101000011000101110001110 ;
        1469: q <= 32'b00111101011101001000110101011100 ;
        1470: q <= 32'b10111100101100010001111101010110 ;
        1471: q <= 32'b00111101000001000100011011001111 ;
        1472: q <= 32'b10111101010111110011100100011111 ;
        1473: q <= 32'b10111100001111001110100010111001 ;
        1474: q <= 32'b00111101100000111010000000101110 ;
        1475: q <= 32'b00111100100110000110100111000111 ;
        1476: q <= 32'b10111101000000111010010100010011 ;
        1477: q <= 32'b00111101011111101100100001001000 ;
        1478: q <= 32'b00111101111100101111110110100010 ;
        1479: q <= 32'b10111101010110000001011010011011 ;
        1480: q <= 32'b10111101101011111111110111100100 ;
        1481: q <= 32'b00111101100101100110010011010101 ;
        1482: q <= 32'b00111101111010000010000000001000 ;
        1483: q <= 32'b10111100111101010101001000001001 ;
        1484: q <= 32'b10111101100110011110010101111110 ;
        1485: q <= 32'b10111101101001010011010000010001 ;
        1486: q <= 32'b10111110000010111111110001110010 ;
        1487: q <= 32'b10111101011110100101001001101011 ;
        1488: q <= 32'b00111101000110110010100100101000 ;
        1489: q <= 32'b10111101010001110111111111010011 ;
        1490: q <= 32'b10111101101111001001100001001110 ;
        1491: q <= 32'b10111101101000000001000001100101 ;
        1492: q <= 32'b10111011101011010000110010110110 ;
        1493: q <= 32'b10111101000000001110110101100010 ;
        1494: q <= 32'b00111101100111101101000110100101 ;
        1495: q <= 32'b10111011100011101101111100100110 ;
        1496: q <= 32'b10111101110110110001001110000010 ;
        1497: q <= 32'b10111101100010111010101100111010 ;
        1498: q <= 32'b00111100011100000011101010011100 ;
        1499: q <= 32'b00111101011100110001011011111101 ;
        1500: q <= 32'b00111101101100111000100100101101 ;
        1501: q <= 32'b00111010000110110011010000010001 ;
        1502: q <= 32'b10111011111011101100011001001011 ;
        1503: q <= 32'b10111100010101011101101111010101 ;
        1504: q <= 32'b10111011100010000110101100000000 ;
        1505: q <= 32'b10111100101010110001111111111111 ;
        1506: q <= 32'b10111101111000111000011101111000 ;
        1507: q <= 32'b00111100111100010101001010000010 ;
        1508: q <= 32'b00111101101001111111111010011110 ;
        1509: q <= 32'b00111100010000000100010100101100 ;
        1510: q <= 32'b00111100101111001000110010110001 ;
        1511: q <= 32'b10111100111010110010001000001111 ;
        1512: q <= 32'b00000000000000000000000000000000 ;
        1513: q <= 32'b00000000000000000000000000000000 ;
        1514: q <= 32'b00000000000000000000000000000000 ;
        1515: q <= 32'b00000000000000000000000000000000 ;
        1516: q <= 32'b00000000000000000000000000000000 ;
        1517: q <= 32'b00000000000000000000000000000000 ;
        1518: q <= 32'b00000000000000000000000000000000 ;
        1519: q <= 32'b00000000000000000000000000000000 ;
        1520: q <= 32'b00000000000000000000000000000000 ;
        1521: q <= 32'b00000000000000000000000000000000 ;
        1522: q <= 32'b00000000000000000000000000000000 ;
        1523: q <= 32'b00000000000000000000000000000000 ;
        1524: q <= 32'b00000000000000000000000000000000 ;
        1525: q <= 32'b00000000000000000000000000000000 ;
        1526: q <= 32'b00000000000000000000000000000000 ;
        1527: q <= 32'b00000000000000000000000000000000 ;
        1528: q <= 32'b00000000000000000000000000000000 ;
        1529: q <= 32'b00000000000000000000000000000000 ;
        1530: q <= 32'b00000000000000000000000000000000 ;
        1531: q <= 32'b00000000000000000000000000000000 ;
        1532: q <= 32'b00000000000000000000000000000000 ;
        1533: q <= 32'b00000000000000000000000000000000 ;
        1534: q <= 32'b00000000000000000000000000000000 ;
        1535: q <= 32'b00000000000000000000000000000000 ;
        1536: q <= 32'b00111101010100111110100110101001 ;
        1537: q <= 32'b00111101010111001100111101001000 ;
        1538: q <= 32'b00111100100100111001011111001011 ;
        1539: q <= 32'b00111100011011110101000111000110 ;
        1540: q <= 32'b10111100011011110110000110011010 ;
        1541: q <= 32'b00111101100001000101000010100111 ;
        1542: q <= 32'b00111101010110010000011011111100 ;
        1543: q <= 32'b10111101011001000001100101110100 ;
        1544: q <= 32'b10111100001000111011100100101001 ;
        1545: q <= 32'b00111101001111001100001110001010 ;
        1546: q <= 32'b10111101011000000101100111111110 ;
        1547: q <= 32'b00111101110001101110010011010110 ;
        1548: q <= 32'b00111100111100011011001111111111 ;
        1549: q <= 32'b00111101011001110001010000100001 ;
        1550: q <= 32'b10111100110101100111111110000011 ;
        1551: q <= 32'b10111101111000001111111110010000 ;
        1552: q <= 32'b00111100111001110111011101101011 ;
        1553: q <= 32'b00111100111000100111011101010001 ;
        1554: q <= 32'b00111100011001001111010010110111 ;
        1555: q <= 32'b10111001001010011001111111011111 ;
        1556: q <= 32'b00111101110111111000001111011111 ;
        1557: q <= 32'b10111101011010111110100010101111 ;
        1558: q <= 32'b10111101101110010110101000111011 ;
        1559: q <= 32'b00111101101010100010011110000101 ;
        1560: q <= 32'b10111101001010010001100111111101 ;
        1561: q <= 32'b10111100001000100001110101101101 ;
        1562: q <= 32'b00111101101101011000000000111011 ;
        1563: q <= 32'b00111011110110100101111000100101 ;
        1564: q <= 32'b00111101100110101010011101101101 ;
        1565: q <= 32'b10111100010001000011000100000011 ;
        1566: q <= 32'b00111100001001000000001110100100 ;
        1567: q <= 32'b00111100101111001110011010000100 ;
        1568: q <= 32'b00111101010110011001001111000100 ;
        1569: q <= 32'b00111101011100000011000111001011 ;
        1570: q <= 32'b00111101101011011001010001101001 ;
        1571: q <= 32'b00111101100001100110001001011001 ;
        1572: q <= 32'b10111101011101101001100000010110 ;
        1573: q <= 32'b10111101000001011000111111101011 ;
        1574: q <= 32'b00111101010100010100100110001111 ;
        1575: q <= 32'b00111101100010000111000111110001 ;
        1576: q <= 32'b00111011101010110011010100010111 ;
        1577: q <= 32'b00111101010010011011101100101000 ;
        1578: q <= 32'b00111100100100100010111110110001 ;
        1579: q <= 32'b00111101001011010010110010101001 ;
        1580: q <= 32'b10111100101100000111011001011110 ;
        1581: q <= 32'b10111101010110010010111101110111 ;
        1582: q <= 32'b00111100100100110001111010000101 ;
        1583: q <= 32'b00111101000100010111110111110101 ;
        1584: q <= 32'b00111101111101110101101111011001 ;
        1585: q <= 32'b10111101010101110101100010000110 ;
        1586: q <= 32'b00111100101110000111001110100010 ;
        1587: q <= 32'b10111101101111101101000100010001 ;
        1588: q <= 32'b00111011100011011101001001100110 ;
        1589: q <= 32'b00111101111111111101001001110100 ;
        1590: q <= 32'b00111101100111001000110000001100 ;
        1591: q <= 32'b10111011110010000010010111111110 ;
        1592: q <= 32'b10111101110100100001110100110100 ;
        1593: q <= 32'b00111100100000111111010101011110 ;
        1594: q <= 32'b10111101100010000000011101101000 ;
        1595: q <= 32'b00111101110010101001101011000000 ;
        1596: q <= 32'b00111101100101101111111000011110 ;
        1597: q <= 32'b00111101001110101110010111010110 ;
        1598: q <= 32'b00111011011111100010111010101110 ;
        1599: q <= 32'b10111100010101011110101111001101 ;
        1600: q <= 32'b10111101101001000010011110001110 ;
        1601: q <= 32'b10111011101110000010011011001011 ;
        1602: q <= 32'b00111101110110010111011001011100 ;
        1603: q <= 32'b00111101110000111111111100100000 ;
        1604: q <= 32'b00111100100010010011100011011010 ;
        1605: q <= 32'b00111101101101001100011010001111 ;
        1606: q <= 32'b00111011110101011101000111010101 ;
        1607: q <= 32'b10111100111001100111001111100101 ;
        1608: q <= 32'b10111101001100110001001100111101 ;
        1609: q <= 32'b10111101101011101110111100110010 ;
        1610: q <= 32'b00111110000000011000101010101100 ;
        1611: q <= 32'b00111101000011010110011001111010 ;
        1612: q <= 32'b00111101111100000101110110010010 ;
        1613: q <= 32'b00111011110001011000110001010011 ;
        1614: q <= 32'b00111101001011110111111000001110 ;
        1615: q <= 32'b00111110000110011001100110000110 ;
        1616: q <= 32'b00111101010100100111101101100100 ;
        1617: q <= 32'b10111101101100110111010100101101 ;
        1618: q <= 32'b10111100011011111111101111101000 ;
        1619: q <= 32'b00111101110011000000001001000000 ;
        1620: q <= 32'b10111101100110001011000001110101 ;
        1621: q <= 32'b00111101111100011111000011110000 ;
        1622: q <= 32'b00111101100001110001100100001011 ;
        1623: q <= 32'b00111100001100100010101010010111 ;
        1624: q <= 32'b10111101010000001111011101000000 ;
        1625: q <= 32'b00111011101101100011010110111010 ;
        1626: q <= 32'b00111101010110000011001111000110 ;
        1627: q <= 32'b00111110001001001101110010010001 ;
        1628: q <= 32'b00111110000101101100001011001011 ;
        1629: q <= 32'b10111011101011011111011111101110 ;
        1630: q <= 32'b10111101010101001110101101111001 ;
        1631: q <= 32'b00111101001111110111000010111010 ;
        1632: q <= 32'b00111101101001110110101110000001 ;
        1633: q <= 32'b00111101000001000011001010100000 ;
        1634: q <= 32'b10111101001110101000011111000011 ;
        1635: q <= 32'b00111101001010011100100101110100 ;
        1636: q <= 32'b10111100110101110101011110001001 ;
        1637: q <= 32'b10111101000000001100110000110110 ;
        1638: q <= 32'b10111101000010111110101010110000 ;
        1639: q <= 32'b00111101101110111110001010011101 ;
        1640: q <= 32'b00000000000000000000000000000000 ;
        1641: q <= 32'b00000000000000000000000000000000 ;
        1642: q <= 32'b00000000000000000000000000000000 ;
        1643: q <= 32'b00000000000000000000000000000000 ;
        1644: q <= 32'b00000000000000000000000000000000 ;
        1645: q <= 32'b00000000000000000000000000000000 ;
        1646: q <= 32'b00000000000000000000000000000000 ;
        1647: q <= 32'b00000000000000000000000000000000 ;
        1648: q <= 32'b00000000000000000000000000000000 ;
        1649: q <= 32'b00000000000000000000000000000000 ;
        1650: q <= 32'b00000000000000000000000000000000 ;
        1651: q <= 32'b00000000000000000000000000000000 ;
        1652: q <= 32'b00000000000000000000000000000000 ;
        1653: q <= 32'b00000000000000000000000000000000 ;
        1654: q <= 32'b00000000000000000000000000000000 ;
        1655: q <= 32'b00000000000000000000000000000000 ;
        1656: q <= 32'b00000000000000000000000000000000 ;
        1657: q <= 32'b00000000000000000000000000000000 ;
        1658: q <= 32'b00000000000000000000000000000000 ;
        1659: q <= 32'b00000000000000000000000000000000 ;
        1660: q <= 32'b00000000000000000000000000000000 ;
        1661: q <= 32'b00000000000000000000000000000000 ;
        1662: q <= 32'b00000000000000000000000000000000 ;
        1663: q <= 32'b00000000000000000000000000000000 ;
        1664: q <= 32'b10111101100011011101010110100101 ;
        1665: q <= 32'b10111101100010100011101010101100 ;
        1666: q <= 32'b10111101110010110000011110110011 ;
        1667: q <= 32'b10111101100100001010001010111100 ;
        1668: q <= 32'b00111101100100001011100001110011 ;
        1669: q <= 32'b00111011110010100100000010011100 ;
        1670: q <= 32'b10111100100111001011000111101010 ;
        1671: q <= 32'b10111101101100010010001110111100 ;
        1672: q <= 32'b00111000011010101000010000011110 ;
        1673: q <= 32'b00111101100001011011010110001001 ;
        1674: q <= 32'b00111101101000111011100111110000 ;
        1675: q <= 32'b00111100000011100000010101111001 ;
        1676: q <= 32'b10111101001010100010111111111111 ;
        1677: q <= 32'b00111100011110001111001011111101 ;
        1678: q <= 32'b10111101100100101011011100010100 ;
        1679: q <= 32'b10111101001010000111101111001110 ;
        1680: q <= 32'b10111101101100110111001011110011 ;
        1681: q <= 32'b10111100011010011001011010101010 ;
        1682: q <= 32'b10111101101101111111010111000001 ;
        1683: q <= 32'b10111101110001000011111011010110 ;
        1684: q <= 32'b10111100010101110101110001110100 ;
        1685: q <= 32'b10111011000001110101010000000001 ;
        1686: q <= 32'b10111101010110110110110110001000 ;
        1687: q <= 32'b00111011101010010110110101001001 ;
        1688: q <= 32'b00111101100110111111111111011100 ;
        1689: q <= 32'b00111101110000011010110000100110 ;
        1690: q <= 32'b00111100011111100110101000101111 ;
        1691: q <= 32'b00111101001011100000011111010011 ;
        1692: q <= 32'b00111101000010110000111010101100 ;
        1693: q <= 32'b00111101100100010101101001110000 ;
        1694: q <= 32'b00111101100011111110011111010001 ;
        1695: q <= 32'b10111101100010111111110100011001 ;
        1696: q <= 32'b10111101101100100110000001000101 ;
        1697: q <= 32'b10111101101010000010111011110110 ;
        1698: q <= 32'b10111101011011111000001101101011 ;
        1699: q <= 32'b10111010101100011001011000011101 ;
        1700: q <= 32'b10111100101010011010110101000110 ;
        1701: q <= 32'b10111101010000010110101110011100 ;
        1702: q <= 32'b00111101010011000001110001100111 ;
        1703: q <= 32'b10111101101100001000000111011100 ;
        1704: q <= 32'b00111100101101110100101111111000 ;
        1705: q <= 32'b00111100111101011110110101111111 ;
        1706: q <= 32'b00111100110001111111110110100010 ;
        1707: q <= 32'b00111100110101001100110100101101 ;
        1708: q <= 32'b10111101101000100010101001001011 ;
        1709: q <= 32'b10111100111111010011100011100110 ;
        1710: q <= 32'b00111100110101001001110011100101 ;
        1711: q <= 32'b00111100100000111000000101010001 ;
        1712: q <= 32'b00111100111100111111100101000111 ;
        1713: q <= 32'b00111101101010000010101100011010 ;
        1714: q <= 32'b00111101000110101001000110111010 ;
        1715: q <= 32'b00111101100001100000100011110011 ;
        1716: q <= 32'b10111110000100001110001000111000 ;
        1717: q <= 32'b10111100100101100100110110010011 ;
        1718: q <= 32'b10111101101010101010101010110000 ;
        1719: q <= 32'b00111101101000001100000010010011 ;
        1720: q <= 32'b00111100101010100110001110111000 ;
        1721: q <= 32'b00111101010100111100000100010011 ;
        1722: q <= 32'b00111100100111001001111000011100 ;
        1723: q <= 32'b10111101101100101100101100110000 ;
        1724: q <= 32'b00111100110100010001110001110010 ;
        1725: q <= 32'b00111100111011011001010000100010 ;
        1726: q <= 32'b10111101101011010101000110010101 ;
        1727: q <= 32'b00111101001101010100100000100110 ;
        1728: q <= 32'b00111100110101110110010000001011 ;
        1729: q <= 32'b00111011101110101010100101101111 ;
        1730: q <= 32'b00111100100000011110011011000010 ;
        1731: q <= 32'b00111100110110111010101111100001 ;
        1732: q <= 32'b10111101101110110000100111001111 ;
        1733: q <= 32'b10111101100010101001011111101011 ;
        1734: q <= 32'b10111101100100100111010010011011 ;
        1735: q <= 32'b00111101101001000110110111111101 ;
        1736: q <= 32'b00111101000111000010000001100110 ;
        1737: q <= 32'b10111101100100001001011100000010 ;
        1738: q <= 32'b00111101000110010100101011000101 ;
        1739: q <= 32'b00111101101000011010010001011101 ;
        1740: q <= 32'b00111101001100001110010000010000 ;
        1741: q <= 32'b00111101101000011100111100001000 ;
        1742: q <= 32'b10111101000101100010001110000101 ;
        1743: q <= 32'b10111101100100110011111110111010 ;
        1744: q <= 32'b00111011010111110110000001001001 ;
        1745: q <= 32'b10111100100110100010110011001011 ;
        1746: q <= 32'b10111100110101010101001110100101 ;
        1747: q <= 32'b10111101011100111010000000011000 ;
        1748: q <= 32'b00111101100111101101000100010000 ;
        1749: q <= 32'b10111100111011101100111110111001 ;
        1750: q <= 32'b00111101100101100001011111010101 ;
        1751: q <= 32'b10111100101011111111111010100010 ;
        1752: q <= 32'b00111101100101011101001100011011 ;
        1753: q <= 32'b00111100100101111111100110011000 ;
        1754: q <= 32'b10111011110110101101111010101111 ;
        1755: q <= 32'b00111101110101010101110110011100 ;
        1756: q <= 32'b10111101100001100000011111101110 ;
        1757: q <= 32'b00111101110010101000011010010100 ;
        1758: q <= 32'b00111101110100010010101010010010 ;
        1759: q <= 32'b10111101010101100111001011000100 ;
        1760: q <= 32'b10111101101101100111111011100011 ;
        1761: q <= 32'b10111101001011100010101111110100 ;
        1762: q <= 32'b10111101101100111011001100000110 ;
        1763: q <= 32'b00111011000000011001010001000010 ;
        1764: q <= 32'b00111100001001111111101101000001 ;
        1765: q <= 32'b00111101100011100111010001010001 ;
        1766: q <= 32'b00111101000101111100100011011100 ;
        1767: q <= 32'b00111101000001111100010101111111 ;
        1768: q <= 32'b00000000000000000000000000000000 ;
        1769: q <= 32'b00000000000000000000000000000000 ;
        1770: q <= 32'b00000000000000000000000000000000 ;
        1771: q <= 32'b00000000000000000000000000000000 ;
        1772: q <= 32'b00000000000000000000000000000000 ;
        1773: q <= 32'b00000000000000000000000000000000 ;
        1774: q <= 32'b00000000000000000000000000000000 ;
        1775: q <= 32'b00000000000000000000000000000000 ;
        1776: q <= 32'b00000000000000000000000000000000 ;
        1777: q <= 32'b00000000000000000000000000000000 ;
        1778: q <= 32'b00000000000000000000000000000000 ;
        1779: q <= 32'b00000000000000000000000000000000 ;
        1780: q <= 32'b00000000000000000000000000000000 ;
        1781: q <= 32'b00000000000000000000000000000000 ;
        1782: q <= 32'b00000000000000000000000000000000 ;
        1783: q <= 32'b00000000000000000000000000000000 ;
        1784: q <= 32'b00000000000000000000000000000000 ;
        1785: q <= 32'b00000000000000000000000000000000 ;
        1786: q <= 32'b00000000000000000000000000000000 ;
        1787: q <= 32'b00000000000000000000000000000000 ;
        1788: q <= 32'b00000000000000000000000000000000 ;
        1789: q <= 32'b00000000000000000000000000000000 ;
        1790: q <= 32'b00000000000000000000000000000000 ;
        1791: q <= 32'b00000000000000000000000000000000 ;
        1792: q <= 32'b10111100111110000111011011111010 ;
        1793: q <= 32'b10111011100001001010011110110111 ;
        1794: q <= 32'b00111011101100111001100110000100 ;
        1795: q <= 32'b10111101001011010101011010101011 ;
        1796: q <= 32'b00111101010011101010000000001011 ;
        1797: q <= 32'b10111101100100000000111101001110 ;
        1798: q <= 32'b00111101000000101110011101001111 ;
        1799: q <= 32'b00111101000101111110100011001101 ;
        1800: q <= 32'b00111100100100001110110110111100 ;
        1801: q <= 32'b00111110000111111110000111001101 ;
        1802: q <= 32'b10111101000111110111111001000010 ;
        1803: q <= 32'b10111100100111110100001001010001 ;
        1804: q <= 32'b10111101011010101100111100110010 ;
        1805: q <= 32'b10111101101000101101100100110100 ;
        1806: q <= 32'b10111100110010010100101000011110 ;
        1807: q <= 32'b10111011011111101111011100011011 ;
        1808: q <= 32'b00111101101000001111111101111111 ;
        1809: q <= 32'b10111110010010110110011101001010 ;
        1810: q <= 32'b10111100000111001010100011000000 ;
        1811: q <= 32'b00111110011101010010100111110111 ;
        1812: q <= 32'b10111100101100010110001111011000 ;
        1813: q <= 32'b00111110000001001111101010100101 ;
        1814: q <= 32'b00111010100011100000011010011001 ;
        1815: q <= 32'b10111110000011110000010011001001 ;
        1816: q <= 32'b00111101000010000101010101010111 ;
        1817: q <= 32'b00111101010101100110110111001101 ;
        1818: q <= 32'b10111101111001101011001000000011 ;
        1819: q <= 32'b00111101100011101001100101101010 ;
        1820: q <= 32'b00111101101001000011000100010011 ;
        1821: q <= 32'b00111101000011011011111011111100 ;
        1822: q <= 32'b00111101110100100101100110101001 ;
        1823: q <= 32'b10111110001111010001110101001110 ;
        1824: q <= 32'b00111101001111101100010010001000 ;
        1825: q <= 32'b00111101101010000010100000010001 ;
        1826: q <= 32'b00111101110011001100110000011110 ;
        1827: q <= 32'b00111100010100001001010001010101 ;
        1828: q <= 32'b10111101111100110000011110010101 ;
        1829: q <= 32'b10111101101101000101101110101011 ;
        1830: q <= 32'b10111101110001101010000010011101 ;
        1831: q <= 32'b10111101110000101101110001010011 ;
        1832: q <= 32'b00111101010100100111001100000100 ;
        1833: q <= 32'b00111100001100001101101111000001 ;
        1834: q <= 32'b10111101001100110110100001001001 ;
        1835: q <= 32'b10111101011111100000000111000011 ;
        1836: q <= 32'b10111101011101001001001100011101 ;
        1837: q <= 32'b00111100101011110101110001001100 ;
        1838: q <= 32'b10111101001000011111101110011000 ;
        1839: q <= 32'b00111101011011110011010011011101 ;
        1840: q <= 32'b10111101100100110101100001100110 ;
        1841: q <= 32'b10111101011110100000000100110010 ;
        1842: q <= 32'b10111101100101101100100101001101 ;
        1843: q <= 32'b10111101100001001111101010101010 ;
        1844: q <= 32'b10111101101110111111000011010010 ;
        1845: q <= 32'b10111011111001111111001111101001 ;
        1846: q <= 32'b00111101100111001111110100110001 ;
        1847: q <= 32'b00111101011110010100101001001101 ;
        1848: q <= 32'b00111100001100010111110000110101 ;
        1849: q <= 32'b10111110001101000011101010000100 ;
        1850: q <= 32'b10111100010111010001100111001101 ;
        1851: q <= 32'b10111101010110010010010011010001 ;
        1852: q <= 32'b10111100001100101011010100000111 ;
        1853: q <= 32'b10111101100000111101001011000110 ;
        1854: q <= 32'b10111110000100000111110111100100 ;
        1855: q <= 32'b10111101010011011011000001001110 ;
        1856: q <= 32'b10111101111001100000111100100111 ;
        1857: q <= 32'b10111110000010100000111111010101 ;
        1858: q <= 32'b00111100111010111100111001111010 ;
        1859: q <= 32'b00111100110110111110011110100110 ;
        1860: q <= 32'b10111100010111001101110010101111 ;
        1861: q <= 32'b10111100010010111001101111010010 ;
        1862: q <= 32'b10111100110111011001111010111001 ;
        1863: q <= 32'b10111100101011000111100101110100 ;
        1864: q <= 32'b00111101011001101101101100011101 ;
        1865: q <= 32'b10111101001011101001101001011101 ;
        1866: q <= 32'b10111110000010101001011101011010 ;
        1867: q <= 32'b10111010111101111000101101110110 ;
        1868: q <= 32'b10111101000111111000110000101111 ;
        1869: q <= 32'b10111101000000100000110110101010 ;
        1870: q <= 32'b10111100001001000001000100100000 ;
        1871: q <= 32'b10111101110011011000100000000101 ;
        1872: q <= 32'b00111101100011000110100100111111 ;
        1873: q <= 32'b00111101101000101010011010110111 ;
        1874: q <= 32'b10111100111011001100000011110100 ;
        1875: q <= 32'b10111110000010001110000011011011 ;
        1876: q <= 32'b00111110000000000100010100111100 ;
        1877: q <= 32'b00111101010111000110101001111111 ;
        1878: q <= 32'b00111100110010101110001111100010 ;
        1879: q <= 32'b10111101000101010100101011011010 ;
        1880: q <= 32'b00111100111011101011011011110010 ;
        1881: q <= 32'b10111101010101000011000000011010 ;
        1882: q <= 32'b10111101101001101011011110110101 ;
        1883: q <= 32'b10111101110011100000111101110011 ;
        1884: q <= 32'b00111101001101110010101001000101 ;
        1885: q <= 32'b10111101000000010110111010001111 ;
        1886: q <= 32'b00111101011000001101100101100010 ;
        1887: q <= 32'b10111101000101110111000010010111 ;
        1888: q <= 32'b00111100101010101001011110101010 ;
        1889: q <= 32'b00111100000110100100100101011000 ;
        1890: q <= 32'b10111100100100111001000110001111 ;
        1891: q <= 32'b10111110000011000001100110111100 ;
        1892: q <= 32'b10111101011100000111111101110011 ;
        1893: q <= 32'b10111011001100110100000000000110 ;
        1894: q <= 32'b00111011000001101100011100111011 ;
        1895: q <= 32'b10111101101011000011011000010110 ;
        1896: q <= 32'b00000000000000000000000000000000 ;
        1897: q <= 32'b00000000000000000000000000000000 ;
        1898: q <= 32'b00000000000000000000000000000000 ;
        1899: q <= 32'b00000000000000000000000000000000 ;
        1900: q <= 32'b00000000000000000000000000000000 ;
        1901: q <= 32'b00000000000000000000000000000000 ;
        1902: q <= 32'b00000000000000000000000000000000 ;
        1903: q <= 32'b00000000000000000000000000000000 ;
        1904: q <= 32'b00000000000000000000000000000000 ;
        1905: q <= 32'b00000000000000000000000000000000 ;
        1906: q <= 32'b00000000000000000000000000000000 ;
        1907: q <= 32'b00000000000000000000000000000000 ;
        1908: q <= 32'b00000000000000000000000000000000 ;
        1909: q <= 32'b00000000000000000000000000000000 ;
        1910: q <= 32'b00000000000000000000000000000000 ;
        1911: q <= 32'b00000000000000000000000000000000 ;
        1912: q <= 32'b00000000000000000000000000000000 ;
        1913: q <= 32'b00000000000000000000000000000000 ;
        1914: q <= 32'b00000000000000000000000000000000 ;
        1915: q <= 32'b00000000000000000000000000000000 ;
        1916: q <= 32'b00000000000000000000000000000000 ;
        1917: q <= 32'b00000000000000000000000000000000 ;
        1918: q <= 32'b00000000000000000000000000000000 ;
        1919: q <= 32'b00000000000000000000000000000000 ;
        1920: q <= 32'b00111101100101100100001110010110 ;
        1921: q <= 32'b00111011000010111011000001100000 ;
        1922: q <= 32'b10111101011101111000001101000100 ;
        1923: q <= 32'b10111101000100110011100000111001 ;
        1924: q <= 32'b10111101111111101101111111010100 ;
        1925: q <= 32'b10111110000010000001011011011010 ;
        1926: q <= 32'b00111100100001011111111111110011 ;
        1927: q <= 32'b10111011111001111111010011111100 ;
        1928: q <= 32'b10111100101100111111111101001100 ;
        1929: q <= 32'b00111101000111101111101001010110 ;
        1930: q <= 32'b10111101111111110000110010011000 ;
        1931: q <= 32'b10111101001110011101000111011101 ;
        1932: q <= 32'b10111101011001101000001001110101 ;
        1933: q <= 32'b00111101100010101000010001100011 ;
        1934: q <= 32'b00111110000010001011111101010111 ;
        1935: q <= 32'b10111101001011100110001011101011 ;
        1936: q <= 32'b10111101100010110010100110111000 ;
        1937: q <= 32'b00111011111110010111101110110000 ;
        1938: q <= 32'b10111101110100011101011001111110 ;
        1939: q <= 32'b10111101011111011111011100001011 ;
        1940: q <= 32'b00111010011110010111000000100111 ;
        1941: q <= 32'b10111101100011010001001001110110 ;
        1942: q <= 32'b10111011001111100100110010011100 ;
        1943: q <= 32'b10111100110000000100111100011001 ;
        1944: q <= 32'b00111100111111110001100101000101 ;
        1945: q <= 32'b00111100011111010111001111101001 ;
        1946: q <= 32'b10111100001110111010011000111001 ;
        1947: q <= 32'b10111100010111011001000011010100 ;
        1948: q <= 32'b00111101101000001001001001110000 ;
        1949: q <= 32'b00111101000010001110101001001000 ;
        1950: q <= 32'b10111100011011011100000101101101 ;
        1951: q <= 32'b00111011000110001000010000111110 ;
        1952: q <= 32'b00111101110101001001011001011010 ;
        1953: q <= 32'b10111100100011110101010011101100 ;
        1954: q <= 32'b10111101001110000100111001101010 ;
        1955: q <= 32'b00111100111100101001010111100010 ;
        1956: q <= 32'b10111110000001011011001001111110 ;
        1957: q <= 32'b10111101010010001000010001000101 ;
        1958: q <= 32'b10111101110101100100001110101001 ;
        1959: q <= 32'b10111100100011101010100000100010 ;
        1960: q <= 32'b00111110001000001100010110111111 ;
        1961: q <= 32'b10111000100010100101001110111011 ;
        1962: q <= 32'b00111110000001101000011101110010 ;
        1963: q <= 32'b10111101100100010111111010001110 ;
        1964: q <= 32'b10111101100111101001001110110011 ;
        1965: q <= 32'b00111101000011110111100111100010 ;
        1966: q <= 32'b10111101010010100010110010111101 ;
        1967: q <= 32'b00111101000001110111000000101010 ;
        1968: q <= 32'b00111100110001011010100010001100 ;
        1969: q <= 32'b10111101101110011111101101001010 ;
        1970: q <= 32'b10111100100001111001001000011101 ;
        1971: q <= 32'b00111101001001011001001001010111 ;
        1972: q <= 32'b00111110001000100000000100100010 ;
        1973: q <= 32'b00111101100011111010001001001010 ;
        1974: q <= 32'b10111101100010111111001010001011 ;
        1975: q <= 32'b10111101101110111101111101101000 ;
        1976: q <= 32'b10111100101000001001110000100011 ;
        1977: q <= 32'b10111100100111101100001100101001 ;
        1978: q <= 32'b00111101111101100100001110010001 ;
        1979: q <= 32'b00111101010100010100111100111100 ;
        1980: q <= 32'b00111101110010100000000010010110 ;
        1981: q <= 32'b10111100111111000110100111010110 ;
        1982: q <= 32'b00111100111010101111000011000011 ;
        1983: q <= 32'b10111101101001011111011010001010 ;
        1984: q <= 32'b10111101100101000000010010100101 ;
        1985: q <= 32'b10111011100110001100110011100110 ;
        1986: q <= 32'b10111100100100110010110100001001 ;
        1987: q <= 32'b10111100010010010011010001100110 ;
        1988: q <= 32'b00111101110111001001100110010110 ;
        1989: q <= 32'b00111100101110000001110110010000 ;
        1990: q <= 32'b10111100010101110001101100101110 ;
        1991: q <= 32'b10111101011100111010011010111011 ;
        1992: q <= 32'b00111101100010001111110110110000 ;
        1993: q <= 32'b10111100100110000000111001110011 ;
        1994: q <= 32'b10111101100010110010001100110111 ;
        1995: q <= 32'b10111101011101010101001000100010 ;
        1996: q <= 32'b10111101100000110000000110100110 ;
        1997: q <= 32'b10111101101000101011000010101101 ;
        1998: q <= 32'b10111101000001111101011110111110 ;
        1999: q <= 32'b10111100110010001001100010010111 ;
        2000: q <= 32'b10111100111111011011100110100010 ;
        2001: q <= 32'b00111110000000100001001110101110 ;
        2002: q <= 32'b10111110000111100001001100010001 ;
        2003: q <= 32'b00111101011001000011110000010110 ;
        2004: q <= 32'b00111101110010011101101110111111 ;
        2005: q <= 32'b10111100101100110001001111011111 ;
        2006: q <= 32'b10111101000001101001011110100001 ;
        2007: q <= 32'b00111011100110100111011000101101 ;
        2008: q <= 32'b10111101000001101000001011100101 ;
        2009: q <= 32'b10111100111100110011001101111001 ;
        2010: q <= 32'b10111011111101101000111011110011 ;
        2011: q <= 32'b10111110000101000001000010000110 ;
        2012: q <= 32'b00111101001010110011111010010110 ;
        2013: q <= 32'b00111100011000000111001010000100 ;
        2014: q <= 32'b00111101000001001100101110001001 ;
        2015: q <= 32'b00111100111110100011111010110010 ;
        2016: q <= 32'b00111100100011010101101011011101 ;
        2017: q <= 32'b00111100110011111101011111111110 ;
        2018: q <= 32'b10111101010111000100010110010011 ;
        2019: q <= 32'b10111100101001111110010010101000 ;
        2020: q <= 32'b00111101000001010100000101001101 ;
        2021: q <= 32'b00111101100000000010110101101000 ;
        2022: q <= 32'b10111101000111001010010010001110 ;
        2023: q <= 32'b10111001100000100010111000010100 ;
        2024: q <= 32'b00000000000000000000000000000000 ;
        2025: q <= 32'b00000000000000000000000000000000 ;
        2026: q <= 32'b00000000000000000000000000000000 ;
        2027: q <= 32'b00000000000000000000000000000000 ;
        2028: q <= 32'b00000000000000000000000000000000 ;
        2029: q <= 32'b00000000000000000000000000000000 ;
        2030: q <= 32'b00000000000000000000000000000000 ;
        2031: q <= 32'b00000000000000000000000000000000 ;
        2032: q <= 32'b00000000000000000000000000000000 ;
        2033: q <= 32'b00000000000000000000000000000000 ;
        2034: q <= 32'b00000000000000000000000000000000 ;
        2035: q <= 32'b00000000000000000000000000000000 ;
        2036: q <= 32'b00000000000000000000000000000000 ;
        2037: q <= 32'b00000000000000000000000000000000 ;
        2038: q <= 32'b00000000000000000000000000000000 ;
        2039: q <= 32'b00000000000000000000000000000000 ;
        2040: q <= 32'b00000000000000000000000000000000 ;
        2041: q <= 32'b00000000000000000000000000000000 ;
        2042: q <= 32'b00000000000000000000000000000000 ;
        2043: q <= 32'b00000000000000000000000000000000 ;
        2044: q <= 32'b00000000000000000000000000000000 ;
        2045: q <= 32'b00000000000000000000000000000000 ;
        2046: q <= 32'b00000000000000000000000000000000 ;
        2047: q <= 32'b00000000000000000000000000000000 ;
        2048: q <= 32'b10111101101101011000001010110100 ;
        2049: q <= 32'b00111100001000101110100000111001 ;
        2050: q <= 32'b00111100110101100001100111000100 ;
        2051: q <= 32'b00111101110001000011111101001001 ;
        2052: q <= 32'b00111100101000111110111001110001 ;
        2053: q <= 32'b10111110001001111101111001111000 ;
        2054: q <= 32'b00111100111111101011110001111010 ;
        2055: q <= 32'b00111101101010100011000101001011 ;
        2056: q <= 32'b10111101101101110001101100011100 ;
        2057: q <= 32'b00111101001010101100100110000011 ;
        2058: q <= 32'b10111101110111001001011100011000 ;
        2059: q <= 32'b10111101100000110000111100100101 ;
        2060: q <= 32'b00111101001010011011011001101111 ;
        2061: q <= 32'b10111110000001101100001101011110 ;
        2062: q <= 32'b00111110000100100110100110110010 ;
        2063: q <= 32'b10111100011001101010001000001100 ;
        2064: q <= 32'b10111101111011111111110011001110 ;
        2065: q <= 32'b10111100000000010010000001110010 ;
        2066: q <= 32'b00111110000001011110010001000110 ;
        2067: q <= 32'b00111101000000001101100001010100 ;
        2068: q <= 32'b10111101100011111101110111100000 ;
        2069: q <= 32'b00111101011110010111000010101110 ;
        2070: q <= 32'b10111101010000100010011000100100 ;
        2071: q <= 32'b00111011100100010100000001101100 ;
        2072: q <= 32'b10111100100101100010111100111001 ;
        2073: q <= 32'b10111100001101111001010110101100 ;
        2074: q <= 32'b00111101010010101111111001100110 ;
        2075: q <= 32'b00111101100101111011001010011010 ;
        2076: q <= 32'b10111101011000101110110010011110 ;
        2077: q <= 32'b10111101110010000101001111001100 ;
        2078: q <= 32'b10111101101000110000001100001110 ;
        2079: q <= 32'b00111100110111010101111100010010 ;
        2080: q <= 32'b00111101000001011111010011001010 ;
        2081: q <= 32'b00111101111001010011000101110100 ;
        2082: q <= 32'b10111100111100001011100001100001 ;
        2083: q <= 32'b10111101000110010001101000111011 ;
        2084: q <= 32'b00111101001011001001110110001111 ;
        2085: q <= 32'b00111011010111111000000110101101 ;
        2086: q <= 32'b00111101100010110101111100110011 ;
        2087: q <= 32'b10111100101110111101111101111111 ;
        2088: q <= 32'b00111101100111111001111100001001 ;
        2089: q <= 32'b10111101011001000101010001101001 ;
        2090: q <= 32'b00111100101011010010111101001110 ;
        2091: q <= 32'b10111101001011100001101010100111 ;
        2092: q <= 32'b10111101101110101011000101111100 ;
        2093: q <= 32'b10111100010001101001000001001100 ;
        2094: q <= 32'b10111100001011100000011101100010 ;
        2095: q <= 32'b00111011100011011001111000011011 ;
        2096: q <= 32'b10111011110011100000100011110000 ;
        2097: q <= 32'b10111101001100101111000110010010 ;
        2098: q <= 32'b10111101100111111100011000100101 ;
        2099: q <= 32'b00111101000101000000000111111101 ;
        2100: q <= 32'b00111101000010111100111000010111 ;
        2101: q <= 32'b10111101100001111001000100111000 ;
        2102: q <= 32'b10111110000001110001010001001001 ;
        2103: q <= 32'b10111101110001001010001010010010 ;
        2104: q <= 32'b10111100110001000001100111111110 ;
        2105: q <= 32'b00111101001111111000010100010111 ;
        2106: q <= 32'b10111101100110110001010001101010 ;
        2107: q <= 32'b10111101010101000011011101000010 ;
        2108: q <= 32'b00111101100000100101110101010011 ;
        2109: q <= 32'b00111100110111000010101011001011 ;
        2110: q <= 32'b10111101111001110010110100110001 ;
        2111: q <= 32'b00111100101001000111101010111001 ;
        2112: q <= 32'b10111100010110100010010001110010 ;
        2113: q <= 32'b00111101101110110000001110001011 ;
        2114: q <= 32'b00111100101111010100010111101101 ;
        2115: q <= 32'b10111100000110101001100110011100 ;
        2116: q <= 32'b10111100110001101110010011101110 ;
        2117: q <= 32'b00111011101001000101000011000101 ;
        2118: q <= 32'b00111100101010110011100110001011 ;
        2119: q <= 32'b10111100001101101000000011000101 ;
        2120: q <= 32'b00111101011100101110001011011000 ;
        2121: q <= 32'b10111101100000110110000101011100 ;
        2122: q <= 32'b00111011001010110010011011001010 ;
        2123: q <= 32'b10111101100100000110110110001110 ;
        2124: q <= 32'b00111101011101100110010100010010 ;
        2125: q <= 32'b00111011100101010101111100110100 ;
        2126: q <= 32'b00111101101001110111011100110001 ;
        2127: q <= 32'b10111011000011111111110111010011 ;
        2128: q <= 32'b10111110000111100010111100010001 ;
        2129: q <= 32'b10111011000011010100011110110100 ;
        2130: q <= 32'b00111100011111101001000000011011 ;
        2131: q <= 32'b10111100111000111111110011001110 ;
        2132: q <= 32'b00111101101000101101101110010001 ;
        2133: q <= 32'b00111101000101110100100001111100 ;
        2134: q <= 32'b00111100101100010001110111000000 ;
        2135: q <= 32'b00111100011100011101100110000000 ;
        2136: q <= 32'b10111101101100011011010110001100 ;
        2137: q <= 32'b00111101011111011001001110001111 ;
        2138: q <= 32'b00111101101110111001111100011001 ;
        2139: q <= 32'b00111101110010001101100100001001 ;
        2140: q <= 32'b10111101010000011110010011001101 ;
        2141: q <= 32'b00111101110010000111111110111110 ;
        2142: q <= 32'b10111101001111100010000101001101 ;
        2143: q <= 32'b00111100100010111101111100000110 ;
        2144: q <= 32'b00111101101001001001001001011101 ;
        2145: q <= 32'b00111101010111110110111101101010 ;
        2146: q <= 32'b00111101101010010000001011010111 ;
        2147: q <= 32'b00111100001011100100111001001011 ;
        2148: q <= 32'b10111100111101001110010111100111 ;
        2149: q <= 32'b00111101011010001100000100001110 ;
        2150: q <= 32'b00111100011101100100000010110101 ;
        2151: q <= 32'b00111010100011001011011010011000 ;
        2152: q <= 32'b00000000000000000000000000000000 ;
        2153: q <= 32'b00000000000000000000000000000000 ;
        2154: q <= 32'b00000000000000000000000000000000 ;
        2155: q <= 32'b00000000000000000000000000000000 ;
        2156: q <= 32'b00000000000000000000000000000000 ;
        2157: q <= 32'b00000000000000000000000000000000 ;
        2158: q <= 32'b00000000000000000000000000000000 ;
        2159: q <= 32'b00000000000000000000000000000000 ;
        2160: q <= 32'b00000000000000000000000000000000 ;
        2161: q <= 32'b00000000000000000000000000000000 ;
        2162: q <= 32'b00000000000000000000000000000000 ;
        2163: q <= 32'b00000000000000000000000000000000 ;
        2164: q <= 32'b00000000000000000000000000000000 ;
        2165: q <= 32'b00000000000000000000000000000000 ;
        2166: q <= 32'b00000000000000000000000000000000 ;
        2167: q <= 32'b00000000000000000000000000000000 ;
        2168: q <= 32'b00000000000000000000000000000000 ;
        2169: q <= 32'b00000000000000000000000000000000 ;
        2170: q <= 32'b00000000000000000000000000000000 ;
        2171: q <= 32'b00000000000000000000000000000000 ;
        2172: q <= 32'b00000000000000000000000000000000 ;
        2173: q <= 32'b00000000000000000000000000000000 ;
        2174: q <= 32'b00000000000000000000000000000000 ;
        2175: q <= 32'b00000000000000000000000000000000 ;
        2176: q <= 32'b10111100100100000011101001110110 ;
        2177: q <= 32'b10111110010011111100000111101010 ;
        2178: q <= 32'b00111101111011101100011011001110 ;
        2179: q <= 32'b00111101111000110001111011011101 ;
        2180: q <= 32'b00111101100101100101000111100101 ;
        2181: q <= 32'b10111100111001110110011000011010 ;
        2182: q <= 32'b10111100110011001110010111000101 ;
        2183: q <= 32'b00111101101000110010011100010011 ;
        2184: q <= 32'b00111101010000001110001000101111 ;
        2185: q <= 32'b10111100000101100101000111010110 ;
        2186: q <= 32'b00111110000001010101010011110000 ;
        2187: q <= 32'b00111101011110000100111011011100 ;
        2188: q <= 32'b00111101101100111011111110000000 ;
        2189: q <= 32'b00111100011010111011101100010001 ;
        2190: q <= 32'b00111101011101101101001110011011 ;
        2191: q <= 32'b10111101101000111101110110011010 ;
        2192: q <= 32'b10111100101111011000111000101010 ;
        2193: q <= 32'b00111100110000001111011100111101 ;
        2194: q <= 32'b00111101110111101011101000000001 ;
        2195: q <= 32'b00111110000001010100001100100010 ;
        2196: q <= 32'b00111100101000111101100001000001 ;
        2197: q <= 32'b10111101001111010100011111100000 ;
        2198: q <= 32'b10111101011000100000110001010011 ;
        2199: q <= 32'b10111011101101110001111010001000 ;
        2200: q <= 32'b00111101100101000111111000101110 ;
        2201: q <= 32'b10111101010101011101110011111101 ;
        2202: q <= 32'b10111101101100010111001001000011 ;
        2203: q <= 32'b10111101110110001100011000111110 ;
        2204: q <= 32'b00111011100001111110100011011101 ;
        2205: q <= 32'b00111110011000010101100010110011 ;
        2206: q <= 32'b00111011001000110000011010111011 ;
        2207: q <= 32'b10111101101001100101011101111011 ;
        2208: q <= 32'b10111100010111111101101000001001 ;
        2209: q <= 32'b10111011110010110110001010101010 ;
        2210: q <= 32'b10111101011001011110110001001000 ;
        2211: q <= 32'b00111101000101110000101110001010 ;
        2212: q <= 32'b00111011101110001110100111110110 ;
        2213: q <= 32'b10111101111100001101001101001111 ;
        2214: q <= 32'b10111101011101000011110011110100 ;
        2215: q <= 32'b00111101100010010001000110000111 ;
        2216: q <= 32'b10111101110110100101100000011110 ;
        2217: q <= 32'b00111101001110001100010111001111 ;
        2218: q <= 32'b00111010011011010110100110100001 ;
        2219: q <= 32'b10111101000000000101100001011111 ;
        2220: q <= 32'b00111101000011001010111100001010 ;
        2221: q <= 32'b00111100101111101110101111110010 ;
        2222: q <= 32'b00111100000000011011011000110000 ;
        2223: q <= 32'b10111011011011000101001100110000 ;
        2224: q <= 32'b00111101010111000000101011101011 ;
        2225: q <= 32'b10111101101000011000101111101011 ;
        2226: q <= 32'b10111101110110011010001001011101 ;
        2227: q <= 32'b00111101011110000001001001101110 ;
        2228: q <= 32'b00111100110001100111001111010110 ;
        2229: q <= 32'b10111100010001010100011111010100 ;
        2230: q <= 32'b00111100010000011100010100110101 ;
        2231: q <= 32'b00111110001000100100110000100101 ;
        2232: q <= 32'b00111110010001110100001001101011 ;
        2233: q <= 32'b00111101101101011010110100010010 ;
        2234: q <= 32'b00111101000100001111111001111111 ;
        2235: q <= 32'b10111101001010010000101111100000 ;
        2236: q <= 32'b10111101001111010001110111001111 ;
        2237: q <= 32'b10111101101001010001000111010010 ;
        2238: q <= 32'b00111101100011001011000111110001 ;
        2239: q <= 32'b10111101110011100101011100101111 ;
        2240: q <= 32'b10111101001011011010110011011100 ;
        2241: q <= 32'b10111101000110001101110110000011 ;
        2242: q <= 32'b10111101111101111001100010101111 ;
        2243: q <= 32'b10111101100011110010100110100111 ;
        2244: q <= 32'b10111100100110000001010101001011 ;
        2245: q <= 32'b00111101100100001101000100000010 ;
        2246: q <= 32'b00111101100100011000110011011110 ;
        2247: q <= 32'b10111110010011010111000100100011 ;
        2248: q <= 32'b10111110000001101001101010101101 ;
        2249: q <= 32'b00111101111101101110000101010110 ;
        2250: q <= 32'b00111101001111001100011011111110 ;
        2251: q <= 32'b00111101100111001011011110000111 ;
        2252: q <= 32'b10111100010110010001011011000101 ;
        2253: q <= 32'b10111101000011001000001010101110 ;
        2254: q <= 32'b00111101100110111000101001101001 ;
        2255: q <= 32'b10111101110101011000111010111001 ;
        2256: q <= 32'b10111101000011010001000011100001 ;
        2257: q <= 32'b00111110001110110111000010111101 ;
        2258: q <= 32'b00111110000111111011000100111010 ;
        2259: q <= 32'b00111110000101011100010101001101 ;
        2260: q <= 32'b00111101101000001111001000111100 ;
        2261: q <= 32'b00111100110001101100110001100001 ;
        2262: q <= 32'b10111101001111011101001111001101 ;
        2263: q <= 32'b00111011111010101110001100101001 ;
        2264: q <= 32'b00111101001011111100000000000011 ;
        2265: q <= 32'b00111101100101100101001000100111 ;
        2266: q <= 32'b00111101110011010111000100000101 ;
        2267: q <= 32'b00111101100111010001011101011011 ;
        2268: q <= 32'b10111101110100100001110010110100 ;
        2269: q <= 32'b00111101100001000100001101010010 ;
        2270: q <= 32'b10111010110010100001011110011110 ;
        2271: q <= 32'b00111011101001001101100100101010 ;
        2272: q <= 32'b00111110010010100011111001111000 ;
        2273: q <= 32'b00111101010011101010000001110100 ;
        2274: q <= 32'b10111101111101110101111001011111 ;
        2275: q <= 32'b00111101110110011001010001101110 ;
        2276: q <= 32'b10111101101000110111010110011000 ;
        2277: q <= 32'b10111100010100110100101011101101 ;
        2278: q <= 32'b00111101110110010001001101001011 ;
        2279: q <= 32'b00111101110101011010001110110011 ;
        2280: q <= 32'b00000000000000000000000000000000 ;
        2281: q <= 32'b00000000000000000000000000000000 ;
        2282: q <= 32'b00000000000000000000000000000000 ;
        2283: q <= 32'b00000000000000000000000000000000 ;
        2284: q <= 32'b00000000000000000000000000000000 ;
        2285: q <= 32'b00000000000000000000000000000000 ;
        2286: q <= 32'b00000000000000000000000000000000 ;
        2287: q <= 32'b00000000000000000000000000000000 ;
        2288: q <= 32'b00000000000000000000000000000000 ;
        2289: q <= 32'b00000000000000000000000000000000 ;
        2290: q <= 32'b00000000000000000000000000000000 ;
        2291: q <= 32'b00000000000000000000000000000000 ;
        2292: q <= 32'b00000000000000000000000000000000 ;
        2293: q <= 32'b00000000000000000000000000000000 ;
        2294: q <= 32'b00000000000000000000000000000000 ;
        2295: q <= 32'b00000000000000000000000000000000 ;
        2296: q <= 32'b00000000000000000000000000000000 ;
        2297: q <= 32'b00000000000000000000000000000000 ;
        2298: q <= 32'b00000000000000000000000000000000 ;
        2299: q <= 32'b00000000000000000000000000000000 ;
        2300: q <= 32'b00000000000000000000000000000000 ;
        2301: q <= 32'b00000000000000000000000000000000 ;
        2302: q <= 32'b00000000000000000000000000000000 ;
        2303: q <= 32'b00000000000000000000000000000000 ;
        2304: q <= 32'b10111101100111011000000100100000 ;
        2305: q <= 32'b00111100111100001001001000111100 ;
        2306: q <= 32'b10111100011001011010000111101111 ;
        2307: q <= 32'b00111110000101001111100111001010 ;
        2308: q <= 32'b10111101101010110010010001001110 ;
        2309: q <= 32'b10111100100100000000100001100101 ;
        2310: q <= 32'b10111110000001111101101111001000 ;
        2311: q <= 32'b00111101011101001011010100111110 ;
        2312: q <= 32'b00111001100111111010001010000001 ;
        2313: q <= 32'b10111101100101111010000000111101 ;
        2314: q <= 32'b00111101100100101001100101111010 ;
        2315: q <= 32'b00111101010001011001001101000111 ;
        2316: q <= 32'b10111100010110110111101011010011 ;
        2317: q <= 32'b10111101000110110110010111000111 ;
        2318: q <= 32'b10111100110010010010101000111010 ;
        2319: q <= 32'b00111110000010101100110000001001 ;
        2320: q <= 32'b10111100001101100110001110000010 ;
        2321: q <= 32'b00111101100010001110001000110100 ;
        2322: q <= 32'b00111101100011101001010110000111 ;
        2323: q <= 32'b10111101110110101000110100110011 ;
        2324: q <= 32'b00111100010010111000010001100000 ;
        2325: q <= 32'b00111101001011000001111011000001 ;
        2326: q <= 32'b00111101100011100111111110000011 ;
        2327: q <= 32'b10111101110100010010110010010101 ;
        2328: q <= 32'b10111101110101111010000111100101 ;
        2329: q <= 32'b00111101010000100100011011111110 ;
        2330: q <= 32'b00111101011011110001001111111111 ;
        2331: q <= 32'b00111101011001001101101100010111 ;
        2332: q <= 32'b10111101100011110000011010100101 ;
        2333: q <= 32'b00111101111100111110001111001000 ;
        2334: q <= 32'b10111101111000001101011010011010 ;
        2335: q <= 32'b10111101111010101101000011100100 ;
        2336: q <= 32'b10111101101010101110100100010100 ;
        2337: q <= 32'b10111010110001010010001001100010 ;
        2338: q <= 32'b00111101100110111111000000100100 ;
        2339: q <= 32'b00111101011111111111110101100100 ;
        2340: q <= 32'b00111101111010101100101101111011 ;
        2341: q <= 32'b10111101000000000011010101000100 ;
        2342: q <= 32'b00111101010101111111001000111111 ;
        2343: q <= 32'b00111101001000000101101111100001 ;
        2344: q <= 32'b00111110001001011101101011100000 ;
        2345: q <= 32'b00111100011111010111000111001001 ;
        2346: q <= 32'b10111100111001101001111001001111 ;
        2347: q <= 32'b10111100111000100111111011011110 ;
        2348: q <= 32'b10111101100110111111111100110000 ;
        2349: q <= 32'b00111010111010111011100011010100 ;
        2350: q <= 32'b00111100001110111111100100000101 ;
        2351: q <= 32'b10111100110110100111010010101111 ;
        2352: q <= 32'b00111100011101111111000111100011 ;
        2353: q <= 32'b00111101110011101001110001000010 ;
        2354: q <= 32'b00111101101101110001101111110111 ;
        2355: q <= 32'b00111101100101011010110010100111 ;
        2356: q <= 32'b10111101001100000010110100011101 ;
        2357: q <= 32'b00111110000001010001111001100000 ;
        2358: q <= 32'b10111101100101100000011001111111 ;
        2359: q <= 32'b00111100110010010100001010011111 ;
        2360: q <= 32'b00111100001111001010000110011001 ;
        2361: q <= 32'b10111110000010100111001000010100 ;
        2362: q <= 32'b10111101000001000100111101000100 ;
        2363: q <= 32'b10111101000001000001011110001011 ;
        2364: q <= 32'b10111100111001100000010001110111 ;
        2365: q <= 32'b10111100001011010100010110011001 ;
        2366: q <= 32'b10111101000101101011000010000100 ;
        2367: q <= 32'b10111101100100011110011101111001 ;
        2368: q <= 32'b10111101111100100100001100010011 ;
        2369: q <= 32'b00111101001110100001111000111001 ;
        2370: q <= 32'b10111101100101001000110001110010 ;
        2371: q <= 32'b10111101010100100101110111110000 ;
        2372: q <= 32'b00111101011111110001011111100010 ;
        2373: q <= 32'b10111100110101010100100110000111 ;
        2374: q <= 32'b10111101001011111010000011010001 ;
        2375: q <= 32'b00111101000110101111001000000010 ;
        2376: q <= 32'b00111101100101000101011000010000 ;
        2377: q <= 32'b10111110000000011000101011001011 ;
        2378: q <= 32'b00111101011110111100001111001100 ;
        2379: q <= 32'b10111100001111000101111110101101 ;
        2380: q <= 32'b10111100011100111100001001010011 ;
        2381: q <= 32'b10111101000000110001011100110010 ;
        2382: q <= 32'b10111101011011100001101000000000 ;
        2383: q <= 32'b10111101100111010010010000010111 ;
        2384: q <= 32'b00111110001100000110001100010111 ;
        2385: q <= 32'b00111110010001011001000101100101 ;
        2386: q <= 32'b00111101011110111011001111111000 ;
        2387: q <= 32'b10111110000101010111011111110111 ;
        2388: q <= 32'b00111101000011001011011000101110 ;
        2389: q <= 32'b10111101101100010111001001001010 ;
        2390: q <= 32'b10111101000000000001011001111101 ;
        2391: q <= 32'b10111101010111010111111100110001 ;
        2392: q <= 32'b10111100110111010000010010011000 ;
        2393: q <= 32'b00111101001101111111011111011111 ;
        2394: q <= 32'b00111101100010110110111101011110 ;
        2395: q <= 32'b10111101001100101110001000001000 ;
        2396: q <= 32'b10111110010010000101001101010001 ;
        2397: q <= 32'b00111101011110011101001100101000 ;
        2398: q <= 32'b10111011100010101001000000011111 ;
        2399: q <= 32'b00111101110110100001010111111101 ;
        2400: q <= 32'b10111101101010111110100110001010 ;
        2401: q <= 32'b00111101101000001010001000010110 ;
        2402: q <= 32'b00111101011110110001010110000001 ;
        2403: q <= 32'b00111101101001001001000110110001 ;
        2404: q <= 32'b10111101000111101110011101011011 ;
        2405: q <= 32'b10111101100101001111110101111001 ;
        2406: q <= 32'b00111101101011010011000110101011 ;
        2407: q <= 32'b10111100001011000011011100010000 ;
        2408: q <= 32'b00000000000000000000000000000000 ;
        2409: q <= 32'b00000000000000000000000000000000 ;
        2410: q <= 32'b00000000000000000000000000000000 ;
        2411: q <= 32'b00000000000000000000000000000000 ;
        2412: q <= 32'b00000000000000000000000000000000 ;
        2413: q <= 32'b00000000000000000000000000000000 ;
        2414: q <= 32'b00000000000000000000000000000000 ;
        2415: q <= 32'b00000000000000000000000000000000 ;
        2416: q <= 32'b00000000000000000000000000000000 ;
        2417: q <= 32'b00000000000000000000000000000000 ;
        2418: q <= 32'b00000000000000000000000000000000 ;
        2419: q <= 32'b00000000000000000000000000000000 ;
        2420: q <= 32'b00000000000000000000000000000000 ;
        2421: q <= 32'b00000000000000000000000000000000 ;
        2422: q <= 32'b00000000000000000000000000000000 ;
        2423: q <= 32'b00000000000000000000000000000000 ;
        2424: q <= 32'b00000000000000000000000000000000 ;
        2425: q <= 32'b00000000000000000000000000000000 ;
        2426: q <= 32'b00000000000000000000000000000000 ;
        2427: q <= 32'b00000000000000000000000000000000 ;
        2428: q <= 32'b00000000000000000000000000000000 ;
        2429: q <= 32'b00000000000000000000000000000000 ;
        2430: q <= 32'b00000000000000000000000000000000 ;
        2431: q <= 32'b00000000000000000000000000000000 ;
        2432: q <= 32'b00111101011111010110100101110110 ;
        2433: q <= 32'b00111011011100011100010101111111 ;
        2434: q <= 32'b10111101010100001111011010110000 ;
        2435: q <= 32'b00111100101001110110111100100011 ;
        2436: q <= 32'b00111101110011110000001010001000 ;
        2437: q <= 32'b00111101110100000110101011100111 ;
        2438: q <= 32'b10111101011111101101000010100110 ;
        2439: q <= 32'b00111100001101011000100001100010 ;
        2440: q <= 32'b00111101101011000010010100011101 ;
        2441: q <= 32'b00111101101110111010011101000110 ;
        2442: q <= 32'b00111100111001010011111000000111 ;
        2443: q <= 32'b10111101111001100101001010010001 ;
        2444: q <= 32'b00111100111011010011101110011101 ;
        2445: q <= 32'b10111101010001110011011110001010 ;
        2446: q <= 32'b10111101001101011000101110011100 ;
        2447: q <= 32'b10111011001111000100010011000100 ;
        2448: q <= 32'b00111101111010011010010011001001 ;
        2449: q <= 32'b00111100010001101110110110010100 ;
        2450: q <= 32'b10111110001000110010111000011101 ;
        2451: q <= 32'b00111101110001111000100000011111 ;
        2452: q <= 32'b00111101100101100101001001101001 ;
        2453: q <= 32'b00111011111101110011101101101100 ;
        2454: q <= 32'b00111101001111101001100100001011 ;
        2455: q <= 32'b10111101110010001101000001110001 ;
        2456: q <= 32'b00111101010001111000001010110101 ;
        2457: q <= 32'b00111011011110010110010010001010 ;
        2458: q <= 32'b00111101001001001111100101100010 ;
        2459: q <= 32'b10111101010101010011111111110011 ;
        2460: q <= 32'b10111011101001000001101100101100 ;
        2461: q <= 32'b10111100011010011001000001011111 ;
        2462: q <= 32'b00111100000001100011001011111011 ;
        2463: q <= 32'b00111101011100111101011010111100 ;
        2464: q <= 32'b10111100110111100111100111001110 ;
        2465: q <= 32'b00111101010101010101110101100111 ;
        2466: q <= 32'b10111100101010100000010000001011 ;
        2467: q <= 32'b00111101110000010111100010110000 ;
        2468: q <= 32'b10111101101110001010000001000111 ;
        2469: q <= 32'b00111101010111001100110110111110 ;
        2470: q <= 32'b00111101101001110011110001111100 ;
        2471: q <= 32'b10111101101111011101101100110111 ;
        2472: q <= 32'b00111010110010011011100111000001 ;
        2473: q <= 32'b10111101010010010101110110010101 ;
        2474: q <= 32'b00111101100111011011111110011010 ;
        2475: q <= 32'b10111101001010110100010001100011 ;
        2476: q <= 32'b10111101111000000110000101110000 ;
        2477: q <= 32'b00111101110011100010110100001000 ;
        2478: q <= 32'b00111101101100111010000001011011 ;
        2479: q <= 32'b10111011001110000110000101011101 ;
        2480: q <= 32'b10111100001100001111100010101100 ;
        2481: q <= 32'b00111100011100100001101100010000 ;
        2482: q <= 32'b00111100110111101100001111011010 ;
        2483: q <= 32'b00111101101010010101111111011111 ;
        2484: q <= 32'b00111101011110101001101110110100 ;
        2485: q <= 32'b10111100000000010110001101110000 ;
        2486: q <= 32'b00111101110000101100110101110010 ;
        2487: q <= 32'b00111101011011010000001100101100 ;
        2488: q <= 32'b00111100101110111000111111001100 ;
        2489: q <= 32'b00111011001000011010111010110110 ;
        2490: q <= 32'b00111110000100011100001111100100 ;
        2491: q <= 32'b10111101100111010001011101101111 ;
        2492: q <= 32'b10111100011111111011001010101100 ;
        2493: q <= 32'b10111100011110111000110001001111 ;
        2494: q <= 32'b00111100101101111001010010101011 ;
        2495: q <= 32'b00111101001111101010100111100111 ;
        2496: q <= 32'b10111101101101000111001000101010 ;
        2497: q <= 32'b10111101111010110111011000110111 ;
        2498: q <= 32'b10111101000000001001100111100100 ;
        2499: q <= 32'b00111101011000001101100111111100 ;
        2500: q <= 32'b00111110000000001010010001000110 ;
        2501: q <= 32'b10111101010110010000111010011100 ;
        2502: q <= 32'b10111101011000100000010010011101 ;
        2503: q <= 32'b00111101001000010110110000101111 ;
        2504: q <= 32'b10111101011110101011111110001000 ;
        2505: q <= 32'b10111011011010111011010000000110 ;
        2506: q <= 32'b10111110000100011101011111001011 ;
        2507: q <= 32'b00111101101100011101100000010100 ;
        2508: q <= 32'b00111101101110110100111001110100 ;
        2509: q <= 32'b10111101011110110010001001011101 ;
        2510: q <= 32'b00111101001101010100101100000011 ;
        2511: q <= 32'b10111100010111111110101001010011 ;
        2512: q <= 32'b00111100111001110100101011100011 ;
        2513: q <= 32'b00111101111101101010010101001100 ;
        2514: q <= 32'b00111100000010010001101110100101 ;
        2515: q <= 32'b10111101110100011011001100011110 ;
        2516: q <= 32'b00111101111110000000101001011110 ;
        2517: q <= 32'b00111101001110110011001100110100 ;
        2518: q <= 32'b10111101111101100111110000000011 ;
        2519: q <= 32'b10111101000110010101111011110100 ;
        2520: q <= 32'b00111101011000000010110000011100 ;
        2521: q <= 32'b00111101000001100100010010111010 ;
        2522: q <= 32'b10111100001001000110010001000111 ;
        2523: q <= 32'b10111110001011110000001001110010 ;
        2524: q <= 32'b00111101110111101110010110110111 ;
        2525: q <= 32'b00111100100101110100110001110100 ;
        2526: q <= 32'b00111101110001000111100011100001 ;
        2527: q <= 32'b10111100111111100110101011100100 ;
        2528: q <= 32'b10111100111100100001001111010010 ;
        2529: q <= 32'b00111100110010111111001010001011 ;
        2530: q <= 32'b10111110000110110101011111011110 ;
        2531: q <= 32'b10111101000110010111011000101000 ;
        2532: q <= 32'b10111101001101010010010111011001 ;
        2533: q <= 32'b10111011101100011001010010110000 ;
        2534: q <= 32'b00111100001110001001100110111010 ;
        2535: q <= 32'b10111100011111010111111101001100 ;
        2536: q <= 32'b00000000000000000000000000000000 ;
        2537: q <= 32'b00000000000000000000000000000000 ;
        2538: q <= 32'b00000000000000000000000000000000 ;
        2539: q <= 32'b00000000000000000000000000000000 ;
        2540: q <= 32'b00000000000000000000000000000000 ;
        2541: q <= 32'b00000000000000000000000000000000 ;
        2542: q <= 32'b00000000000000000000000000000000 ;
        2543: q <= 32'b00000000000000000000000000000000 ;
        2544: q <= 32'b00000000000000000000000000000000 ;
        2545: q <= 32'b00000000000000000000000000000000 ;
        2546: q <= 32'b00000000000000000000000000000000 ;
        2547: q <= 32'b00000000000000000000000000000000 ;
        2548: q <= 32'b00000000000000000000000000000000 ;
        2549: q <= 32'b00000000000000000000000000000000 ;
        2550: q <= 32'b00000000000000000000000000000000 ;
        2551: q <= 32'b00000000000000000000000000000000 ;
        2552: q <= 32'b00000000000000000000000000000000 ;
        2553: q <= 32'b00000000000000000000000000000000 ;
        2554: q <= 32'b00000000000000000000000000000000 ;
        2555: q <= 32'b00000000000000000000000000000000 ;
        2556: q <= 32'b00000000000000000000000000000000 ;
        2557: q <= 32'b00000000000000000000000000000000 ;
        2558: q <= 32'b00000000000000000000000000000000 ;
        2559: q <= 32'b00000000000000000000000000000000 ;
        2560: q <= 32'b00111101100001111110011000110010 ;
        2561: q <= 32'b10111100000001001010101010111000 ;
        2562: q <= 32'b10111101000100000111000101000111 ;
        2563: q <= 32'b00111101010111001100100010100100 ;
        2564: q <= 32'b10111101011001100010011011011001 ;
        2565: q <= 32'b10111100000000011111111110010110 ;
        2566: q <= 32'b00111101011101000110011010100111 ;
        2567: q <= 32'b10111110000111111110001000000110 ;
        2568: q <= 32'b00111101110110001100100100010111 ;
        2569: q <= 32'b00111101101011011001110111100110 ;
        2570: q <= 32'b10111101100110001001000101000010 ;
        2571: q <= 32'b10111101100001000001111111000001 ;
        2572: q <= 32'b00111101011101000100001101001010 ;
        2573: q <= 32'b10111100101010101100001100110011 ;
        2574: q <= 32'b00111011110000110100100101001001 ;
        2575: q <= 32'b00111110010011000011111001000101 ;
        2576: q <= 32'b10111100011100111001011001110111 ;
        2577: q <= 32'b00111100100101100100111100000011 ;
        2578: q <= 32'b00111101000000010011010100010000 ;
        2579: q <= 32'b00111100101010000101100100001110 ;
        2580: q <= 32'b00111101011010000001001100101100 ;
        2581: q <= 32'b00111100000000100101111111111010 ;
        2582: q <= 32'b00111101010101010111000000001110 ;
        2583: q <= 32'b10111100101011010110100000111100 ;
        2584: q <= 32'b10111110001010010101011100100101 ;
        2585: q <= 32'b00111100010101101101100011110011 ;
        2586: q <= 32'b00111101010101011101110001111111 ;
        2587: q <= 32'b10111101100011111010100000101001 ;
        2588: q <= 32'b10111100001101110101000111001001 ;
        2589: q <= 32'b00111101011001100011010101010111 ;
        2590: q <= 32'b10111101111111011100100011100000 ;
        2591: q <= 32'b00111101110101100100001010010100 ;
        2592: q <= 32'b00111101100101011111001000000011 ;
        2593: q <= 32'b10111100010110110101010001010110 ;
        2594: q <= 32'b00111110000011001101100010100110 ;
        2595: q <= 32'b10111100010101110010110001000100 ;
        2596: q <= 32'b10111101111000111110111110100011 ;
        2597: q <= 32'b00111101110010101011100011111001 ;
        2598: q <= 32'b00111101000000001001011011010101 ;
        2599: q <= 32'b10111100000000011001001110100000 ;
        2600: q <= 32'b00111101110001000101100000011100 ;
        2601: q <= 32'b00111101101110101111110100110100 ;
        2602: q <= 32'b00111101101111010100011111111100 ;
        2603: q <= 32'b10111100111111111110011011011101 ;
        2604: q <= 32'b00111101100000110111100011100000 ;
        2605: q <= 32'b00111010100011011110010010111101 ;
        2606: q <= 32'b10111101010101010101110001000100 ;
        2607: q <= 32'b10111011100111111000111111111001 ;
        2608: q <= 32'b10111100110110101001101101101000 ;
        2609: q <= 32'b10111101000101010001110111001110 ;
        2610: q <= 32'b00111100111100101001010100000111 ;
        2611: q <= 32'b10111011000110011110110001001100 ;
        2612: q <= 32'b10111101100010101101110111010110 ;
        2613: q <= 32'b10111101010100110011110011011111 ;
        2614: q <= 32'b10111110000000000001111000011111 ;
        2615: q <= 32'b10111101010000111100100010000011 ;
        2616: q <= 32'b10111011110011111110101011001110 ;
        2617: q <= 32'b00111100111000101000000001010101 ;
        2618: q <= 32'b00111100011010011111111001100001 ;
        2619: q <= 32'b10111110000001111101011101100110 ;
        2620: q <= 32'b00111101111110011010011011010100 ;
        2621: q <= 32'b10111100111101000100100100100001 ;
        2622: q <= 32'b00111011111100000010110100111001 ;
        2623: q <= 32'b00111101001011101100001011010100 ;
        2624: q <= 32'b00111010101100011000000110110001 ;
        2625: q <= 32'b10111100101000101011001101001010 ;
        2626: q <= 32'b10111101010110001101011100111111 ;
        2627: q <= 32'b10111101100011111011001000000010 ;
        2628: q <= 32'b00111100110011100011000000011010 ;
        2629: q <= 32'b10111101010100101000000011000100 ;
        2630: q <= 32'b10111011100111100000111111101010 ;
        2631: q <= 32'b00111100111010101000110111101100 ;
        2632: q <= 32'b10111100001111001110010100000000 ;
        2633: q <= 32'b10111100001111110101000011111110 ;
        2634: q <= 32'b00111101001101101111011001011011 ;
        2635: q <= 32'b00111101100011000101101011010101 ;
        2636: q <= 32'b10111101010110010001011001110011 ;
        2637: q <= 32'b10111011010101110110110010101010 ;
        2638: q <= 32'b10111101001011111000001101111010 ;
        2639: q <= 32'b10111101110110011011000001101100 ;
        2640: q <= 32'b10111110000011110011010101000000 ;
        2641: q <= 32'b10111011101010110110001011110000 ;
        2642: q <= 32'b10111101111101010001011110010001 ;
        2643: q <= 32'b00111101011010110110010111001010 ;
        2644: q <= 32'b00111101101100010001101100101101 ;
        2645: q <= 32'b10111101000101011001101100101000 ;
        2646: q <= 32'b00111101010101011101110100101010 ;
        2647: q <= 32'b10111101000010000011101011100011 ;
        2648: q <= 32'b10111110000001111010010111100101 ;
        2649: q <= 32'b10111101010101011000110101010011 ;
        2650: q <= 32'b00111100100000101101100010110000 ;
        2651: q <= 32'b10111110001001101110110001001000 ;
        2652: q <= 32'b10111110000100000111011011101110 ;
        2653: q <= 32'b00111010000000010101011110100000 ;
        2654: q <= 32'b10111101000111110100100111000101 ;
        2655: q <= 32'b10111101001100100010111001010000 ;
        2656: q <= 32'b10111101000010010010110000010001 ;
        2657: q <= 32'b10111101100000000011010001010000 ;
        2658: q <= 32'b00111100101100001110111111111011 ;
        2659: q <= 32'b10111101101110100101001010100010 ;
        2660: q <= 32'b00111100110110010100101011100101 ;
        2661: q <= 32'b10111101011011001101110110010110 ;
        2662: q <= 32'b00111101101001001101010011111111 ;
        2663: q <= 32'b10111100111011100001000101000001 ;
        2664: q <= 32'b00000000000000000000000000000000 ;
        2665: q <= 32'b00000000000000000000000000000000 ;
        2666: q <= 32'b00000000000000000000000000000000 ;
        2667: q <= 32'b00000000000000000000000000000000 ;
        2668: q <= 32'b00000000000000000000000000000000 ;
        2669: q <= 32'b00000000000000000000000000000000 ;
        2670: q <= 32'b00000000000000000000000000000000 ;
        2671: q <= 32'b00000000000000000000000000000000 ;
        2672: q <= 32'b00000000000000000000000000000000 ;
        2673: q <= 32'b00000000000000000000000000000000 ;
        2674: q <= 32'b00000000000000000000000000000000 ;
        2675: q <= 32'b00000000000000000000000000000000 ;
        2676: q <= 32'b00000000000000000000000000000000 ;
        2677: q <= 32'b00000000000000000000000000000000 ;
        2678: q <= 32'b00000000000000000000000000000000 ;
        2679: q <= 32'b00000000000000000000000000000000 ;
        2680: q <= 32'b00000000000000000000000000000000 ;
        2681: q <= 32'b00000000000000000000000000000000 ;
        2682: q <= 32'b00000000000000000000000000000000 ;
        2683: q <= 32'b00000000000000000000000000000000 ;
        2684: q <= 32'b00000000000000000000000000000000 ;
        2685: q <= 32'b00000000000000000000000000000000 ;
        2686: q <= 32'b00000000000000000000000000000000 ;
        2687: q <= 32'b00000000000000000000000000000000 ;
        2688: q <= 32'b10111011000000010100011101111101 ;
        2689: q <= 32'b00111101100111101100100111110000 ;
        2690: q <= 32'b10111100000100110011100101010001 ;
        2691: q <= 32'b10111101010011011101100100110100 ;
        2692: q <= 32'b00111101100100000011011111010110 ;
        2693: q <= 32'b10111010111010011011101100001100 ;
        2694: q <= 32'b10111101011100100110001001111111 ;
        2695: q <= 32'b10111101001100111000000111010000 ;
        2696: q <= 32'b10111100110110101100011001010101 ;
        2697: q <= 32'b10111101100110010010101110000101 ;
        2698: q <= 32'b00111101101000001010010110010011 ;
        2699: q <= 32'b10111101101101011101111001011001 ;
        2700: q <= 32'b00111101010011100111011101111000 ;
        2701: q <= 32'b00111101101011001101110000101110 ;
        2702: q <= 32'b10111100100100011111111001011100 ;
        2703: q <= 32'b10111101110111000001110001111101 ;
        2704: q <= 32'b10111101010110011000101001000110 ;
        2705: q <= 32'b00111101000110011011111011110000 ;
        2706: q <= 32'b00111101000111000101101111111111 ;
        2707: q <= 32'b00111101001000000000010101000001 ;
        2708: q <= 32'b10111100011010110000001110111011 ;
        2709: q <= 32'b10111100001101011010101111101101 ;
        2710: q <= 32'b00111101110011000101111011110000 ;
        2711: q <= 32'b00111101000111111001001010000101 ;
        2712: q <= 32'b10111101001100100011011111000001 ;
        2713: q <= 32'b10111101101011010000100001011100 ;
        2714: q <= 32'b10111101110010001001100100110111 ;
        2715: q <= 32'b00111101110111010110100111001101 ;
        2716: q <= 32'b10111101110101011001101010111101 ;
        2717: q <= 32'b10111101100000101100101101010010 ;
        2718: q <= 32'b10111101110010000001011100101110 ;
        2719: q <= 32'b00111101000000011100001001011000 ;
        2720: q <= 32'b00111100010101110000010101011110 ;
        2721: q <= 32'b10111011010001000010001001110100 ;
        2722: q <= 32'b10111101001100010101001110011110 ;
        2723: q <= 32'b10111101111011010010011011010001 ;
        2724: q <= 32'b00111101100101001001100111000110 ;
        2725: q <= 32'b00111100111110101001100111101111 ;
        2726: q <= 32'b00111101101001001010101111100100 ;
        2727: q <= 32'b00111100000000110001000011010110 ;
        2728: q <= 32'b10111101010101100111111100101011 ;
        2729: q <= 32'b00111101010101000110000111110100 ;
        2730: q <= 32'b00111101111000110110011001000101 ;
        2731: q <= 32'b10111011000101111110000100100001 ;
        2732: q <= 32'b10111101011010011000100010100010 ;
        2733: q <= 32'b10111100101101110011010001001110 ;
        2734: q <= 32'b00111101101000111101011000110111 ;
        2735: q <= 32'b00111101001101100110110111110100 ;
        2736: q <= 32'b00111101111111000001100011111100 ;
        2737: q <= 32'b00111101000110101111011110111100 ;
        2738: q <= 32'b10111101110010100000110001100011 ;
        2739: q <= 32'b00111101100101010111001101010000 ;
        2740: q <= 32'b00111100001111000010100111001011 ;
        2741: q <= 32'b10111101101011101100000011101111 ;
        2742: q <= 32'b10111110001111101101101101111101 ;
        2743: q <= 32'b10111101100101101101001100000010 ;
        2744: q <= 32'b10111101110100011101111001111000 ;
        2745: q <= 32'b00111101000000011000111100000111 ;
        2746: q <= 32'b00111100011100001001101111111111 ;
        2747: q <= 32'b00111101100010000001101001000110 ;
        2748: q <= 32'b00111101100110000010000101010000 ;
        2749: q <= 32'b10111101110001111111001011110101 ;
        2750: q <= 32'b00111011010101100011001111101010 ;
        2751: q <= 32'b10111011110110011010110111001010 ;
        2752: q <= 32'b10111101011111101110001000100001 ;
        2753: q <= 32'b00111101110010110111000011000001 ;
        2754: q <= 32'b10111101110001101001000110100011 ;
        2755: q <= 32'b00111101101101010001000110010010 ;
        2756: q <= 32'b00111100110110101010110010001001 ;
        2757: q <= 32'b10111101001100101110101100010100 ;
        2758: q <= 32'b00111101111110001011101100000111 ;
        2759: q <= 32'b00111101100011000001111000101101 ;
        2760: q <= 32'b10111101001011110000111011000111 ;
        2761: q <= 32'b00111110000010010111100111100001 ;
        2762: q <= 32'b00111100101100011000010011100111 ;
        2763: q <= 32'b00111101000000010101100000010110 ;
        2764: q <= 32'b00111011001110101001010111111110 ;
        2765: q <= 32'b00111100100011010011010101001010 ;
        2766: q <= 32'b10111011101010011010111001011110 ;
        2767: q <= 32'b10111110001101111101010010000000 ;
        2768: q <= 32'b00111101000011101111110010100000 ;
        2769: q <= 32'b10111101110101011110100111010111 ;
        2770: q <= 32'b10111101011101001001010000101111 ;
        2771: q <= 32'b10111011110101010101111110000001 ;
        2772: q <= 32'b10111100101001111100101101001011 ;
        2773: q <= 32'b00111100111111111111001111110010 ;
        2774: q <= 32'b10111101000110101000001010010010 ;
        2775: q <= 32'b00111100111000001111001011000110 ;
        2776: q <= 32'b10111101001010111100000100011100 ;
        2777: q <= 32'b00111101011001011101111101110011 ;
        2778: q <= 32'b00111101111000000010000001110000 ;
        2779: q <= 32'b00111101111001100110010010100111 ;
        2780: q <= 32'b10111011110100100000000001111011 ;
        2781: q <= 32'b00111101110110011110010011001100 ;
        2782: q <= 32'b10111100101010110011000110011010 ;
        2783: q <= 32'b00111101110000110000001011010001 ;
        2784: q <= 32'b00111100111110100001110000110000 ;
        2785: q <= 32'b00111101100100001111000111111000 ;
        2786: q <= 32'b00111101001010100010110100110110 ;
        2787: q <= 32'b00111101110010101001110011111011 ;
        2788: q <= 32'b00111101100000100010001000000100 ;
        2789: q <= 32'b00111011111000111001001110110011 ;
        2790: q <= 32'b10111101100101010011100010001101 ;
        2791: q <= 32'b10111101100110101101010111100011 ;
        2792: q <= 32'b00000000000000000000000000000000 ;
        2793: q <= 32'b00000000000000000000000000000000 ;
        2794: q <= 32'b00000000000000000000000000000000 ;
        2795: q <= 32'b00000000000000000000000000000000 ;
        2796: q <= 32'b00000000000000000000000000000000 ;
        2797: q <= 32'b00000000000000000000000000000000 ;
        2798: q <= 32'b00000000000000000000000000000000 ;
        2799: q <= 32'b00000000000000000000000000000000 ;
        2800: q <= 32'b00000000000000000000000000000000 ;
        2801: q <= 32'b00000000000000000000000000000000 ;
        2802: q <= 32'b00000000000000000000000000000000 ;
        2803: q <= 32'b00000000000000000000000000000000 ;
        2804: q <= 32'b00000000000000000000000000000000 ;
        2805: q <= 32'b00000000000000000000000000000000 ;
        2806: q <= 32'b00000000000000000000000000000000 ;
        2807: q <= 32'b00000000000000000000000000000000 ;
        2808: q <= 32'b00000000000000000000000000000000 ;
        2809: q <= 32'b00000000000000000000000000000000 ;
        2810: q <= 32'b00000000000000000000000000000000 ;
        2811: q <= 32'b00000000000000000000000000000000 ;
        2812: q <= 32'b00000000000000000000000000000000 ;
        2813: q <= 32'b00000000000000000000000000000000 ;
        2814: q <= 32'b00000000000000000000000000000000 ;
        2815: q <= 32'b00000000000000000000000000000000 ;
        2816: q <= 32'b00111101100101111100001011010111 ;
        2817: q <= 32'b00111101110010100100100001100111 ;
        2818: q <= 32'b10111011010100000010001100010010 ;
        2819: q <= 32'b00111100101110110011010110011110 ;
        2820: q <= 32'b00111100101010011110000011010010 ;
        2821: q <= 32'b00111101001101010101111011100001 ;
        2822: q <= 32'b10111101101011110111011000100001 ;
        2823: q <= 32'b10111101111110110011010101100100 ;
        2824: q <= 32'b10111100001101000001101000111101 ;
        2825: q <= 32'b10111110000011100110010100100110 ;
        2826: q <= 32'b00111011011011000110011000011011 ;
        2827: q <= 32'b10111101100000111010000111010101 ;
        2828: q <= 32'b10111010001010001100100101001101 ;
        2829: q <= 32'b10111100111001110110100000111110 ;
        2830: q <= 32'b10111100101101010000111010111100 ;
        2831: q <= 32'b00111011101000110101110100111101 ;
        2832: q <= 32'b00111101111000101010000110111111 ;
        2833: q <= 32'b00111101000010101011010010111111 ;
        2834: q <= 32'b10111101001101010001010101100011 ;
        2835: q <= 32'b00111101011000011001001111011101 ;
        2836: q <= 32'b00111101000010011111111010100011 ;
        2837: q <= 32'b10111101110101111101100111101111 ;
        2838: q <= 32'b10111100000101100000010100010010 ;
        2839: q <= 32'b10111100110001000101100001100010 ;
        2840: q <= 32'b00111011100010000000011010101010 ;
        2841: q <= 32'b00111100100000010100000000010011 ;
        2842: q <= 32'b10111011101000100110010111010110 ;
        2843: q <= 32'b00111101101100110111010010011100 ;
        2844: q <= 32'b10111101101011110001111110111100 ;
        2845: q <= 32'b00111101110000101011001100110001 ;
        2846: q <= 32'b00111101101111100001011010101110 ;
        2847: q <= 32'b00111101010101101010100000110000 ;
        2848: q <= 32'b10111101110000111000101111110110 ;
        2849: q <= 32'b00111101111010101000011010110011 ;
        2850: q <= 32'b00111100010100111111001100101101 ;
        2851: q <= 32'b10111101000100111100100011100111 ;
        2852: q <= 32'b00111101001001010001001011000110 ;
        2853: q <= 32'b10111011010000101111100000111100 ;
        2854: q <= 32'b10111101011100111100100000100010 ;
        2855: q <= 32'b00111101001000100100100100110000 ;
        2856: q <= 32'b00111100011001011001000101010011 ;
        2857: q <= 32'b10111101011001011011011011010101 ;
        2858: q <= 32'b10111101100010010101111111000011 ;
        2859: q <= 32'b00111100110100111111110110101011 ;
        2860: q <= 32'b10111110000011110100000110001011 ;
        2861: q <= 32'b10111100100001000111010100111111 ;
        2862: q <= 32'b00111101111101011110101010011010 ;
        2863: q <= 32'b10111101010010101110001111000101 ;
        2864: q <= 32'b00111101110100010110101101001101 ;
        2865: q <= 32'b00111100100101001001011110101100 ;
        2866: q <= 32'b10111100010110010110100010000100 ;
        2867: q <= 32'b00111101110001111101101001100111 ;
        2868: q <= 32'b00111101100000111101010000111011 ;
        2869: q <= 32'b00111101010011101011101101111011 ;
        2870: q <= 32'b00111101110101011010100001011110 ;
        2871: q <= 32'b10111101001110011001010011000011 ;
        2872: q <= 32'b00111101010000001111011001100000 ;
        2873: q <= 32'b00111100001100000001111011101000 ;
        2874: q <= 32'b00111011100110000101000000000101 ;
        2875: q <= 32'b10111101001110100110010000100001 ;
        2876: q <= 32'b10111101111100011000011101000011 ;
        2877: q <= 32'b00111100000111011001010110011000 ;
        2878: q <= 32'b00111101111001000010010010010100 ;
        2879: q <= 32'b00111100000100000111000001001000 ;
        2880: q <= 32'b00111101100100010001011111110101 ;
        2881: q <= 32'b10111110010000110100001110000011 ;
        2882: q <= 32'b00111101000011010101100100010101 ;
        2883: q <= 32'b00111101111011011011110111100000 ;
        2884: q <= 32'b10111101110111011101110001111110 ;
        2885: q <= 32'b00111100110010010100011111010010 ;
        2886: q <= 32'b10111011101010100001010111011100 ;
        2887: q <= 32'b00111101000101000101010000100011 ;
        2888: q <= 32'b10111101111011110011100000011010 ;
        2889: q <= 32'b10111101010111111011110001010110 ;
        2890: q <= 32'b10111101001100001101011010101001 ;
        2891: q <= 32'b10111101010100111101011001011001 ;
        2892: q <= 32'b10111101100111101110100010011101 ;
        2893: q <= 32'b00111101100111110011111100010100 ;
        2894: q <= 32'b10111101101001100000011111111011 ;
        2895: q <= 32'b00111101101100011010100001011011 ;
        2896: q <= 32'b10111101001110111000110011000101 ;
        2897: q <= 32'b10111110000100100111100101101000 ;
        2898: q <= 32'b00111110001101111001111111011000 ;
        2899: q <= 32'b00111101111011010100011100010010 ;
        2900: q <= 32'b10111101111100110100001001001110 ;
        2901: q <= 32'b00111101100111100110010100110111 ;
        2902: q <= 32'b10111100100110110110100110000101 ;
        2903: q <= 32'b10111011111011110001110101110110 ;
        2904: q <= 32'b00111101101010001101001101010101 ;
        2905: q <= 32'b00111101010100010010100011101111 ;
        2906: q <= 32'b10111101101101001000010100000101 ;
        2907: q <= 32'b00111101101010101010110110011011 ;
        2908: q <= 32'b10111101011110010111010011110101 ;
        2909: q <= 32'b00111101000011010101111011110000 ;
        2910: q <= 32'b10111100110001011110010001000010 ;
        2911: q <= 32'b00111110000001111000010101001111 ;
        2912: q <= 32'b10111101100110010010001001111001 ;
        2913: q <= 32'b10111100111000110000100100111001 ;
        2914: q <= 32'b00111101111100001110111110101001 ;
        2915: q <= 32'b10111011010110110000110001001011 ;
        2916: q <= 32'b10111100110101010011100000110111 ;
        2917: q <= 32'b10111010111100110101110011010001 ;
        2918: q <= 32'b10111101010010110001001000110110 ;
        2919: q <= 32'b00111100000111000010010011011000 ;
        2920: q <= 32'b00000000000000000000000000000000 ;
        2921: q <= 32'b00000000000000000000000000000000 ;
        2922: q <= 32'b00000000000000000000000000000000 ;
        2923: q <= 32'b00000000000000000000000000000000 ;
        2924: q <= 32'b00000000000000000000000000000000 ;
        2925: q <= 32'b00000000000000000000000000000000 ;
        2926: q <= 32'b00000000000000000000000000000000 ;
        2927: q <= 32'b00000000000000000000000000000000 ;
        2928: q <= 32'b00000000000000000000000000000000 ;
        2929: q <= 32'b00000000000000000000000000000000 ;
        2930: q <= 32'b00000000000000000000000000000000 ;
        2931: q <= 32'b00000000000000000000000000000000 ;
        2932: q <= 32'b00000000000000000000000000000000 ;
        2933: q <= 32'b00000000000000000000000000000000 ;
        2934: q <= 32'b00000000000000000000000000000000 ;
        2935: q <= 32'b00000000000000000000000000000000 ;
        2936: q <= 32'b00000000000000000000000000000000 ;
        2937: q <= 32'b00000000000000000000000000000000 ;
        2938: q <= 32'b00000000000000000000000000000000 ;
        2939: q <= 32'b00000000000000000000000000000000 ;
        2940: q <= 32'b00000000000000000000000000000000 ;
        2941: q <= 32'b00000000000000000000000000000000 ;
        2942: q <= 32'b00000000000000000000000000000000 ;
        2943: q <= 32'b00000000000000000000000000000000 ;
        2944: q <= 32'b00111101100000111110110000010100 ;
        2945: q <= 32'b10111101100110010110011111001010 ;
        2946: q <= 32'b00111100000111101011001010100011 ;
        2947: q <= 32'b00111110000000101100001111101101 ;
        2948: q <= 32'b10111101011110110100111000101011 ;
        2949: q <= 32'b00111101011100010001100101001010 ;
        2950: q <= 32'b00111101100111101111000110001000 ;
        2951: q <= 32'b00111101101011101100001001110111 ;
        2952: q <= 32'b10111100000101001111000110000101 ;
        2953: q <= 32'b10111101110010111010111111000001 ;
        2954: q <= 32'b00111100011100100010100001101101 ;
        2955: q <= 32'b00111011110100111000010001001001 ;
        2956: q <= 32'b00111101011010000001010101111110 ;
        2957: q <= 32'b10111101000111101100111011010011 ;
        2958: q <= 32'b00111101100001100001100010111110 ;
        2959: q <= 32'b00111101011011011110011001000001 ;
        2960: q <= 32'b00111101011111101001011110111001 ;
        2961: q <= 32'b00111100101111101011100110010011 ;
        2962: q <= 32'b00111100111110010101101010101011 ;
        2963: q <= 32'b00111101110011110100110100110101 ;
        2964: q <= 32'b10111101010010000111011010010110 ;
        2965: q <= 32'b10111101111011101001111100000100 ;
        2966: q <= 32'b00111101010100110110100000001010 ;
        2967: q <= 32'b10111011111101111111001111001001 ;
        2968: q <= 32'b00111101100100010110100000001010 ;
        2969: q <= 32'b10111101000011010010001000010100 ;
        2970: q <= 32'b00111101010101111101011000100001 ;
        2971: q <= 32'b10111101101101100111101011101101 ;
        2972: q <= 32'b10111100000100010101000111010011 ;
        2973: q <= 32'b00111101010011010000000001110011 ;
        2974: q <= 32'b10111101101100011110011111010000 ;
        2975: q <= 32'b00111101100111101011111011010000 ;
        2976: q <= 32'b00111101111100001001011011100000 ;
        2977: q <= 32'b00111011110001000111000010100011 ;
        2978: q <= 32'b10111101011010000110000110001100 ;
        2979: q <= 32'b00111101011011101010110110111010 ;
        2980: q <= 32'b00111100101100011001110100101010 ;
        2981: q <= 32'b10111100110010110001000011110001 ;
        2982: q <= 32'b10111100111100111101011010001101 ;
        2983: q <= 32'b10111101100011111010010100000101 ;
        2984: q <= 32'b10111101001111111110111111001010 ;
        2985: q <= 32'b00111101101110000110101000101101 ;
        2986: q <= 32'b10111100100110000111100101110000 ;
        2987: q <= 32'b10111101000110110101001011000110 ;
        2988: q <= 32'b10111101100000111011011111110001 ;
        2989: q <= 32'b00111101000111011010100101011011 ;
        2990: q <= 32'b10111101101010110110001111111001 ;
        2991: q <= 32'b00111101010100110110001111100011 ;
        2992: q <= 32'b10111101100001000000110011011000 ;
        2993: q <= 32'b10111100100111110100101111000010 ;
        2994: q <= 32'b10111101101011010101001010010110 ;
        2995: q <= 32'b00111101100101010011111001001110 ;
        2996: q <= 32'b00111101111110110000110100000000 ;
        2997: q <= 32'b10111101001001110100101001110101 ;
        2998: q <= 32'b00111101010111001110111110000111 ;
        2999: q <= 32'b00111101001011110111011101110011 ;
        3000: q <= 32'b10111001111110101010001010100110 ;
        3001: q <= 32'b00111101110111000000101010101011 ;
        3002: q <= 32'b00111101100100110000101000010100 ;
        3003: q <= 32'b10111101101110101111001011110010 ;
        3004: q <= 32'b10111101110100110011111000101111 ;
        3005: q <= 32'b10111101001010001100000111011111 ;
        3006: q <= 32'b10111010100000110111001101001001 ;
        3007: q <= 32'b00111101101010110000010111010110 ;
        3008: q <= 32'b10111101101110101001101010101011 ;
        3009: q <= 32'b10111101001100100000000010011011 ;
        3010: q <= 32'b10111010110111101110010101000111 ;
        3011: q <= 32'b00111100111111001101111111010000 ;
        3012: q <= 32'b10111101100101001101000111001111 ;
        3013: q <= 32'b10111100101111010010110001100010 ;
        3014: q <= 32'b00111101100100100100011100111000 ;
        3015: q <= 32'b00111100100110010100111110010110 ;
        3016: q <= 32'b10111101000011011100111110011111 ;
        3017: q <= 32'b00111100000000011100100001011000 ;
        3018: q <= 32'b10111100000110100111100111100111 ;
        3019: q <= 32'b10111101010011111011001111010100 ;
        3020: q <= 32'b10111101010101000011011001111111 ;
        3021: q <= 32'b00111100111110101001100100010111 ;
        3022: q <= 32'b10111101010010011011000111110000 ;
        3023: q <= 32'b00111101011100111101010100001111 ;
        3024: q <= 32'b00111101100101110110001010111010 ;
        3025: q <= 32'b10111101100100001010101010001100 ;
        3026: q <= 32'b00111101000111101101000010101001 ;
        3027: q <= 32'b10111101000000001111010111010100 ;
        3028: q <= 32'b00111100100010011101000100001100 ;
        3029: q <= 32'b00111100010100101111101010110100 ;
        3030: q <= 32'b10111101011011000110010010111000 ;
        3031: q <= 32'b10111101100100100011111000111110 ;
        3032: q <= 32'b00111101001101101011110000101100 ;
        3033: q <= 32'b00111101100100000000110000001100 ;
        3034: q <= 32'b10111101010000010110110000110011 ;
        3035: q <= 32'b10111101101101000110110001000111 ;
        3036: q <= 32'b00111101001011111110111000000111 ;
        3037: q <= 32'b10111101101000110111101111000000 ;
        3038: q <= 32'b00111101010000011100111011111001 ;
        3039: q <= 32'b00111101111001000011001100010010 ;
        3040: q <= 32'b10111101010100111000111001001001 ;
        3041: q <= 32'b00111101000110010000100000001001 ;
        3042: q <= 32'b00111101101001000101001100100011 ;
        3043: q <= 32'b00111100111111010010100011011000 ;
        3044: q <= 32'b10111100101101010101001101100001 ;
        3045: q <= 32'b10111100100001010100111111111010 ;
        3046: q <= 32'b00111101001010011101000101010010 ;
        3047: q <= 32'b00111101101001111001001011000010 ;
        3048: q <= 32'b00000000000000000000000000000000 ;
        3049: q <= 32'b00000000000000000000000000000000 ;
        3050: q <= 32'b00000000000000000000000000000000 ;
        3051: q <= 32'b00000000000000000000000000000000 ;
        3052: q <= 32'b00000000000000000000000000000000 ;
        3053: q <= 32'b00000000000000000000000000000000 ;
        3054: q <= 32'b00000000000000000000000000000000 ;
        3055: q <= 32'b00000000000000000000000000000000 ;
        3056: q <= 32'b00000000000000000000000000000000 ;
        3057: q <= 32'b00000000000000000000000000000000 ;
        3058: q <= 32'b00000000000000000000000000000000 ;
        3059: q <= 32'b00000000000000000000000000000000 ;
        3060: q <= 32'b00000000000000000000000000000000 ;
        3061: q <= 32'b00000000000000000000000000000000 ;
        3062: q <= 32'b00000000000000000000000000000000 ;
        3063: q <= 32'b00000000000000000000000000000000 ;
        3064: q <= 32'b00000000000000000000000000000000 ;
        3065: q <= 32'b00000000000000000000000000000000 ;
        3066: q <= 32'b00000000000000000000000000000000 ;
        3067: q <= 32'b00000000000000000000000000000000 ;
        3068: q <= 32'b00000000000000000000000000000000 ;
        3069: q <= 32'b00000000000000000000000000000000 ;
        3070: q <= 32'b00000000000000000000000000000000 ;
        3071: q <= 32'b00000000000000000000000000000000 ;
        3072: q <= 32'b00111100000000011011000011010101 ;
        3073: q <= 32'b10111101010101000101001101010010 ;
        3074: q <= 32'b10111101001010101110100010101110 ;
        3075: q <= 32'b00111100010000101101111011011100 ;
        3076: q <= 32'b10111101011111000000010110100110 ;
        3077: q <= 32'b10111101001010100101101000001000 ;
        3078: q <= 32'b00111101111110000110110110111101 ;
        3079: q <= 32'b10111100111011101011010100100001 ;
        3080: q <= 32'b10111101100100000100110101000110 ;
        3081: q <= 32'b10111011110101011000111010100000 ;
        3082: q <= 32'b00111100110100110010001110001100 ;
        3083: q <= 32'b00111100011111010110101111010011 ;
        3084: q <= 32'b00111100000011100010100001100110 ;
        3085: q <= 32'b00111100101100110001001000010101 ;
        3086: q <= 32'b00111100110111110111110001010000 ;
        3087: q <= 32'b10111101010100100010111100100110 ;
        3088: q <= 32'b10111101110100111010100110100000 ;
        3089: q <= 32'b10111101010111000000110111111111 ;
        3090: q <= 32'b10111101011110100110011111111100 ;
        3091: q <= 32'b00111100011000110010001100101110 ;
        3092: q <= 32'b10111011110001010110010001011110 ;
        3093: q <= 32'b10111100111111100011101010100000 ;
        3094: q <= 32'b00111011000101010000001110011011 ;
        3095: q <= 32'b00111100101110001100110101101011 ;
        3096: q <= 32'b00111100100100011111100100010010 ;
        3097: q <= 32'b10111100101000101110101001101010 ;
        3098: q <= 32'b10111101101100100011111100010101 ;
        3099: q <= 32'b00111011010110011110111001001011 ;
        3100: q <= 32'b10111101000111001000111101011100 ;
        3101: q <= 32'b10111101011101010110100001001100 ;
        3102: q <= 32'b10111100010101101001011011111100 ;
        3103: q <= 32'b10111101011111101100011100001000 ;
        3104: q <= 32'b00111100100001100111110010001001 ;
        3105: q <= 32'b00111100101000111010111111000111 ;
        3106: q <= 32'b10111101001100001011110000010011 ;
        3107: q <= 32'b10111101001011100010101001000011 ;
        3108: q <= 32'b10111101100110000100001000010100 ;
        3109: q <= 32'b00111100111000110100100100110001 ;
        3110: q <= 32'b10111011001010001010011010110100 ;
        3111: q <= 32'b10111101001110001101001001111111 ;
        3112: q <= 32'b10111101001101110100000011100110 ;
        3113: q <= 32'b10111100011000111100111010111011 ;
        3114: q <= 32'b00111101100110001000011011001110 ;
        3115: q <= 32'b00111010111101001101001100110000 ;
        3116: q <= 32'b10111100100100100110110111010001 ;
        3117: q <= 32'b00111101100000101111110011100010 ;
        3118: q <= 32'b10111101000101111000101101110110 ;
        3119: q <= 32'b00111110000111011100110111011000 ;
        3120: q <= 32'b10111101011111100110011000111111 ;
        3121: q <= 32'b10111101101101011101011000001001 ;
        3122: q <= 32'b10111100101011001010111110101001 ;
        3123: q <= 32'b10111100111111100011100110110010 ;
        3124: q <= 32'b10111110000101110100101100111100 ;
        3125: q <= 32'b10111100110001111111100011001111 ;
        3126: q <= 32'b00111101101010011010001100001011 ;
        3127: q <= 32'b10111101101000100011011100010101 ;
        3128: q <= 32'b10111001011101111110011111101101 ;
        3129: q <= 32'b00111011100001111111101001011101 ;
        3130: q <= 32'b00111101011101100100000110011001 ;
        3131: q <= 32'b00111101100110011100100011010111 ;
        3132: q <= 32'b10111100100001110100000011101110 ;
        3133: q <= 32'b10111100111111000101000010011001 ;
        3134: q <= 32'b00111100100100101100011110100111 ;
        3135: q <= 32'b00111100100011100100010100000000 ;
        3136: q <= 32'b00111101110101011001011011001111 ;
        3137: q <= 32'b10111110000110000011101111111010 ;
        3138: q <= 32'b00111101101001001010001000001111 ;
        3139: q <= 32'b00111110000101010100111001110110 ;
        3140: q <= 32'b00111100010010010010111111110111 ;
        3141: q <= 32'b00111100110101111010010111001111 ;
        3142: q <= 32'b10111011000000101110111111000000 ;
        3143: q <= 32'b00111101001010000100011000011010 ;
        3144: q <= 32'b00111101000000011011100001100011 ;
        3145: q <= 32'b10111100100011010001000001011100 ;
        3146: q <= 32'b10111101100111001001011101101011 ;
        3147: q <= 32'b10111101110010100001111010100100 ;
        3148: q <= 32'b10111101001000101011101101100100 ;
        3149: q <= 32'b00111101100111100100001011101100 ;
        3150: q <= 32'b10111101011010010010011100101010 ;
        3151: q <= 32'b00111011010100110011110010000110 ;
        3152: q <= 32'b00111101110001110100011011110001 ;
        3153: q <= 32'b00111101011011111010100101000011 ;
        3154: q <= 32'b10111101110111101011010100110010 ;
        3155: q <= 32'b10111110001111100001001110100110 ;
        3156: q <= 32'b00111101000001010001000111101110 ;
        3157: q <= 32'b10111101000110110100001011000110 ;
        3158: q <= 32'b10111011010001011001101001111000 ;
        3159: q <= 32'b10111101111101011011000111101000 ;
        3160: q <= 32'b10111101101011100010001100010101 ;
        3161: q <= 32'b00111101000100101101010011010000 ;
        3162: q <= 32'b10111100000011000011000100101100 ;
        3163: q <= 32'b10111101100110000111001001001001 ;
        3164: q <= 32'b00111110001101110110011000101110 ;
        3165: q <= 32'b10111100010001011111101000010000 ;
        3166: q <= 32'b00111100111011001100111111010110 ;
        3167: q <= 32'b00111101101011011110100010101101 ;
        3168: q <= 32'b10111110001010001101111110000010 ;
        3169: q <= 32'b00111101010100110111001110110110 ;
        3170: q <= 32'b10111011100000101010011011000101 ;
        3171: q <= 32'b10111100101110000011010010110000 ;
        3172: q <= 32'b00111101100110111011001001001000 ;
        3173: q <= 32'b10111011100011110011000101110001 ;
        3174: q <= 32'b00111101000010101010010110010010 ;
        3175: q <= 32'b00111100001010111100010110111111 ;
        3176: q <= 32'b00000000000000000000000000000000 ;
        3177: q <= 32'b00000000000000000000000000000000 ;
        3178: q <= 32'b00000000000000000000000000000000 ;
        3179: q <= 32'b00000000000000000000000000000000 ;
        3180: q <= 32'b00000000000000000000000000000000 ;
        3181: q <= 32'b00000000000000000000000000000000 ;
        3182: q <= 32'b00000000000000000000000000000000 ;
        3183: q <= 32'b00000000000000000000000000000000 ;
        3184: q <= 32'b00000000000000000000000000000000 ;
        3185: q <= 32'b00000000000000000000000000000000 ;
        3186: q <= 32'b00000000000000000000000000000000 ;
        3187: q <= 32'b00000000000000000000000000000000 ;
        3188: q <= 32'b00000000000000000000000000000000 ;
        3189: q <= 32'b00000000000000000000000000000000 ;
        3190: q <= 32'b00000000000000000000000000000000 ;
        3191: q <= 32'b00000000000000000000000000000000 ;
        3192: q <= 32'b00000000000000000000000000000000 ;
        3193: q <= 32'b00000000000000000000000000000000 ;
        3194: q <= 32'b00000000000000000000000000000000 ;
        3195: q <= 32'b00000000000000000000000000000000 ;
        3196: q <= 32'b00000000000000000000000000000000 ;
        3197: q <= 32'b00000000000000000000000000000000 ;
        3198: q <= 32'b00000000000000000000000000000000 ;
        3199: q <= 32'b00000000000000000000000000000000 ;
        3200: q <= 32'b10111101111110010001110110000100 ;
        3201: q <= 32'b00111101011100011001100101100011 ;
        3202: q <= 32'b00111101010000011101111001000110 ;
        3203: q <= 32'b00111101101000001110110001111001 ;
        3204: q <= 32'b10111000101111010011001000001101 ;
        3205: q <= 32'b00111100101000110011010001100000 ;
        3206: q <= 32'b10111100101111100111001110010010 ;
        3207: q <= 32'b00111101100101100000111010001000 ;
        3208: q <= 32'b10111101011110011000100000101001 ;
        3209: q <= 32'b10111101101111111010010001110110 ;
        3210: q <= 32'b00111101100110111000111110010100 ;
        3211: q <= 32'b00111100110001010000101101110101 ;
        3212: q <= 32'b10111011110111101110111101011011 ;
        3213: q <= 32'b00111101110001000111100111111011 ;
        3214: q <= 32'b00111101001110010000100001000110 ;
        3215: q <= 32'b10111100010001010110000001001000 ;
        3216: q <= 32'b10111101001010110001001101001011 ;
        3217: q <= 32'b00111101110110110000110010110001 ;
        3218: q <= 32'b00111101001010111111110101000000 ;
        3219: q <= 32'b10111100101111001001010000111111 ;
        3220: q <= 32'b10111101111001010010011011100110 ;
        3221: q <= 32'b00111100110100101110111011000011 ;
        3222: q <= 32'b10111100111101011100011001011101 ;
        3223: q <= 32'b00111101000010011001111010000101 ;
        3224: q <= 32'b00111101100101101111010110101111 ;
        3225: q <= 32'b00111101010100100001001000010011 ;
        3226: q <= 32'b10111100111101010011000100101001 ;
        3227: q <= 32'b10111101101101001111110001001010 ;
        3228: q <= 32'b10111011111001001011001010010010 ;
        3229: q <= 32'b00111101111100000111110111111101 ;
        3230: q <= 32'b00111100101110111001100101011101 ;
        3231: q <= 32'b00111101100001001001000000111110 ;
        3232: q <= 32'b10111101010000100011001110101000 ;
        3233: q <= 32'b10111101001001100110001101110000 ;
        3234: q <= 32'b00111100010000111110101001111000 ;
        3235: q <= 32'b10111101110010111010100110110110 ;
        3236: q <= 32'b00111100100101000001100101110011 ;
        3237: q <= 32'b00111101001111000000000110010001 ;
        3238: q <= 32'b00111101100000011100110011110010 ;
        3239: q <= 32'b10111100101001001000001000001001 ;
        3240: q <= 32'b10111101010011100011001010101111 ;
        3241: q <= 32'b10111101011111001011100000010000 ;
        3242: q <= 32'b10111110010010110100000000101000 ;
        3243: q <= 32'b00111100110010011111001011110010 ;
        3244: q <= 32'b00111100001001010010110101101010 ;
        3245: q <= 32'b10111101010010000101000001100011 ;
        3246: q <= 32'b10111101000000011001010100011011 ;
        3247: q <= 32'b10111100000010111100111101110000 ;
        3248: q <= 32'b00111100010000101010100111101100 ;
        3249: q <= 32'b10111100010000000001110100110000 ;
        3250: q <= 32'b00111101011000001011001011011011 ;
        3251: q <= 32'b10111101000111001101001011000000 ;
        3252: q <= 32'b00111101101011011110001000010111 ;
        3253: q <= 32'b10111101101110001001000100111000 ;
        3254: q <= 32'b10111101011010101100101100010100 ;
        3255: q <= 32'b10111101001111100001100100010011 ;
        3256: q <= 32'b10111101001101011101010101011111 ;
        3257: q <= 32'b00111101100101100101001001010101 ;
        3258: q <= 32'b10111101101111011000001111101111 ;
        3259: q <= 32'b00111101100001010000100100010000 ;
        3260: q <= 32'b00111100000101101010100111011111 ;
        3261: q <= 32'b00111100111010001010001101110111 ;
        3262: q <= 32'b00111101100010001111001010100001 ;
        3263: q <= 32'b00111101000110001100011000100011 ;
        3264: q <= 32'b00111101100101010001111010100011 ;
        3265: q <= 32'b00111100000111001110011000111001 ;
        3266: q <= 32'b00111101101010000110111100111000 ;
        3267: q <= 32'b10111011111001101001110000110110 ;
        3268: q <= 32'b10111101101100000011011010111001 ;
        3269: q <= 32'b00111101000101000101001001101010 ;
        3270: q <= 32'b00111101100010011001100000110000 ;
        3271: q <= 32'b10111101001101101001011010111010 ;
        3272: q <= 32'b00111101010101000110001111011111 ;
        3273: q <= 32'b10111100101011100011111001011111 ;
        3274: q <= 32'b00111101100010101100101000100000 ;
        3275: q <= 32'b10111101010101100100101011010101 ;
        3276: q <= 32'b10111101111011011100100111101010 ;
        3277: q <= 32'b10111101100101010100000110011011 ;
        3278: q <= 32'b10111101110000010000101111011000 ;
        3279: q <= 32'b10111101000111000000001110101110 ;
        3280: q <= 32'b10111100011111010110110110111111 ;
        3281: q <= 32'b10111101000111010001110011111101 ;
        3282: q <= 32'b00111110001011000011011001010010 ;
        3283: q <= 32'b00111101000010101111001010100101 ;
        3284: q <= 32'b10111101100100111010010100010100 ;
        3285: q <= 32'b00111101011101011111100010011110 ;
        3286: q <= 32'b00111101110111110111100101100111 ;
        3287: q <= 32'b00111110000001101111011101010111 ;
        3288: q <= 32'b00111101101100100001110111000110 ;
        3289: q <= 32'b00111101010101101110101011101000 ;
        3290: q <= 32'b00111101000110100100010010100111 ;
        3291: q <= 32'b00111101110010011100100111000010 ;
        3292: q <= 32'b00111101010001001111100110010111 ;
        3293: q <= 32'b10111100000110001101001100110010 ;
        3294: q <= 32'b00111101000011111011100011101010 ;
        3295: q <= 32'b00110111110101001111011001111101 ;
        3296: q <= 32'b10111100111100010111100111010000 ;
        3297: q <= 32'b00111101100001100011111110001111 ;
        3298: q <= 32'b10111100011001101000101010100110 ;
        3299: q <= 32'b00111100111101100001001111100000 ;
        3300: q <= 32'b10111101011111010100101011011110 ;
        3301: q <= 32'b10111100100011011111110000011111 ;
        3302: q <= 32'b10111100101001000011100110111000 ;
        3303: q <= 32'b00111101001110110000010000010011 ;
        3304: q <= 32'b00000000000000000000000000000000 ;
        3305: q <= 32'b00000000000000000000000000000000 ;
        3306: q <= 32'b00000000000000000000000000000000 ;
        3307: q <= 32'b00000000000000000000000000000000 ;
        3308: q <= 32'b00000000000000000000000000000000 ;
        3309: q <= 32'b00000000000000000000000000000000 ;
        3310: q <= 32'b00000000000000000000000000000000 ;
        3311: q <= 32'b00000000000000000000000000000000 ;
        3312: q <= 32'b00000000000000000000000000000000 ;
        3313: q <= 32'b00000000000000000000000000000000 ;
        3314: q <= 32'b00000000000000000000000000000000 ;
        3315: q <= 32'b00000000000000000000000000000000 ;
        3316: q <= 32'b00000000000000000000000000000000 ;
        3317: q <= 32'b00000000000000000000000000000000 ;
        3318: q <= 32'b00000000000000000000000000000000 ;
        3319: q <= 32'b00000000000000000000000000000000 ;
        3320: q <= 32'b00000000000000000000000000000000 ;
        3321: q <= 32'b00000000000000000000000000000000 ;
        3322: q <= 32'b00000000000000000000000000000000 ;
        3323: q <= 32'b00000000000000000000000000000000 ;
        3324: q <= 32'b00000000000000000000000000000000 ;
        3325: q <= 32'b00000000000000000000000000000000 ;
        3326: q <= 32'b00000000000000000000000000000000 ;
        3327: q <= 32'b00000000000000000000000000000000 ;
        3328: q <= 32'b00111101010011111110011100100110 ;
        3329: q <= 32'b00111101101111010101101110010010 ;
        3330: q <= 32'b10111100110001100000111100101010 ;
        3331: q <= 32'b10111110001101101101100111110101 ;
        3332: q <= 32'b00111110000110001100111000111011 ;
        3333: q <= 32'b00111110000111110000110001001101 ;
        3334: q <= 32'b10111101110000110100110001111000 ;
        3335: q <= 32'b10111101101011000101110000111011 ;
        3336: q <= 32'b00111101001011100000000001101111 ;
        3337: q <= 32'b00111101100011101101101111011011 ;
        3338: q <= 32'b00111100010100100011001100100010 ;
        3339: q <= 32'b00111101101101111100101101000000 ;
        3340: q <= 32'b10111101001001001100010100100011 ;
        3341: q <= 32'b10111101010101101000001101110101 ;
        3342: q <= 32'b10111101110000110101100001100111 ;
        3343: q <= 32'b10111101100000011001101101100000 ;
        3344: q <= 32'b00111110000010110010100000011111 ;
        3345: q <= 32'b00111100101110010001001000010000 ;
        3346: q <= 32'b00111101101000001011110111101001 ;
        3347: q <= 32'b00111100010011010000110101001101 ;
        3348: q <= 32'b10111001101011011010011100011100 ;
        3349: q <= 32'b00111110000010101000000001101001 ;
        3350: q <= 32'b10111101100000011101101011010111 ;
        3351: q <= 32'b10111100110000011001111010011000 ;
        3352: q <= 32'b10111011101010001111111101010011 ;
        3353: q <= 32'b10111101100001100001100011101011 ;
        3354: q <= 32'b10111110000010011011010011101100 ;
        3355: q <= 32'b00111101110011000011110001110110 ;
        3356: q <= 32'b00111100111110110111100001100110 ;
        3357: q <= 32'b10111110010000100001000101110010 ;
        3358: q <= 32'b00111110000011011110110001110000 ;
        3359: q <= 32'b00111101011100010110011000010111 ;
        3360: q <= 32'b10111101111010100111110001000010 ;
        3361: q <= 32'b00111101011000010111101001001001 ;
        3362: q <= 32'b10111100111000101111011111101111 ;
        3363: q <= 32'b10111101100101011001111101110000 ;
        3364: q <= 32'b00111100100010011001000110000111 ;
        3365: q <= 32'b00111100111100000110000010010011 ;
        3366: q <= 32'b00111101101001110011010000011111 ;
        3367: q <= 32'b10111100110010100111001011000001 ;
        3368: q <= 32'b10111101001001000110000100110010 ;
        3369: q <= 32'b10111100111000100111001111011111 ;
        3370: q <= 32'b00111101111000111111111010100000 ;
        3371: q <= 32'b10111101100001101100100010000000 ;
        3372: q <= 32'b00111100000001010110011101000101 ;
        3373: q <= 32'b00111100011101111111100101110000 ;
        3374: q <= 32'b10111101100110110111100100011111 ;
        3375: q <= 32'b00111101101011010111101111011100 ;
        3376: q <= 32'b00111100100010100011011000010111 ;
        3377: q <= 32'b00111101001000110111010010111010 ;
        3378: q <= 32'b10111100100011001001011100001001 ;
        3379: q <= 32'b00111100110011011011100011011010 ;
        3380: q <= 32'b00111011100001101110000001111011 ;
        3381: q <= 32'b10111101010101101110100011100001 ;
        3382: q <= 32'b00111100011011001000010110101000 ;
        3383: q <= 32'b10111110000001100001011110101000 ;
        3384: q <= 32'b00111110001011011110100000111000 ;
        3385: q <= 32'b00111101101011110100110110000000 ;
        3386: q <= 32'b10111101101011111111110000101011 ;
        3387: q <= 32'b10111101100010010001000110010011 ;
        3388: q <= 32'b00111101000010101110101011001110 ;
        3389: q <= 32'b10111101010010001100001101101011 ;
        3390: q <= 32'b10111101100111110010000101111111 ;
        3391: q <= 32'b10111101001000001100001010110110 ;
        3392: q <= 32'b10111100011100111100001100000011 ;
        3393: q <= 32'b10111100101100101001111000110001 ;
        3394: q <= 32'b10111101000001000111001010100101 ;
        3395: q <= 32'b00111101110000101001001101000000 ;
        3396: q <= 32'b00111100110011110001010000101111 ;
        3397: q <= 32'b10111101100000110000100111110101 ;
        3398: q <= 32'b10111110000000100001110111110010 ;
        3399: q <= 32'b00111101001011001001110101100011 ;
        3400: q <= 32'b00111101101101011111100011010110 ;
        3401: q <= 32'b10111101101000110111000111100000 ;
        3402: q <= 32'b10111101000110010010101101101011 ;
        3403: q <= 32'b00111101000001011111100010001001 ;
        3404: q <= 32'b10111101010110111111101010000101 ;
        3405: q <= 32'b00111101000101101110011000010110 ;
        3406: q <= 32'b10111100001100110101001111101010 ;
        3407: q <= 32'b00111101110010001110100011101011 ;
        3408: q <= 32'b00111101100101001111010000000100 ;
        3409: q <= 32'b10111101000011001000111101101100 ;
        3410: q <= 32'b00111110010101000101000101110000 ;
        3411: q <= 32'b00111110001011100101011000010100 ;
        3412: q <= 32'b00111100101110011101100111001010 ;
        3413: q <= 32'b00111101100110001101111001101100 ;
        3414: q <= 32'b10111101000011001101100110001101 ;
        3415: q <= 32'b10111101100110101010011010110111 ;
        3416: q <= 32'b00111100000000110111011011000010 ;
        3417: q <= 32'b00111011110110000010011010010110 ;
        3418: q <= 32'b10111101101001110100001101111001 ;
        3419: q <= 32'b00111100110001001111010100101010 ;
        3420: q <= 32'b00111101000111110101111100111001 ;
        3421: q <= 32'b00111101101100100101000110100101 ;
        3422: q <= 32'b00111101110001001010010011011011 ;
        3423: q <= 32'b00111100100001011010101110001010 ;
        3424: q <= 32'b00111101010001111011110100110111 ;
        3425: q <= 32'b10111101011110000011001101011101 ;
        3426: q <= 32'b00111110000000110110101010000000 ;
        3427: q <= 32'b00111100001001001010011100110100 ;
        3428: q <= 32'b00111100101100110110010000100110 ;
        3429: q <= 32'b00111101000000111000000111100011 ;
        3430: q <= 32'b00111101010000110011001101001010 ;
        3431: q <= 32'b00111101111001010110100110100100 ;
        3432: q <= 32'b00000000000000000000000000000000 ;
        3433: q <= 32'b00000000000000000000000000000000 ;
        3434: q <= 32'b00000000000000000000000000000000 ;
        3435: q <= 32'b00000000000000000000000000000000 ;
        3436: q <= 32'b00000000000000000000000000000000 ;
        3437: q <= 32'b00000000000000000000000000000000 ;
        3438: q <= 32'b00000000000000000000000000000000 ;
        3439: q <= 32'b00000000000000000000000000000000 ;
        3440: q <= 32'b00000000000000000000000000000000 ;
        3441: q <= 32'b00000000000000000000000000000000 ;
        3442: q <= 32'b00000000000000000000000000000000 ;
        3443: q <= 32'b00000000000000000000000000000000 ;
        3444: q <= 32'b00000000000000000000000000000000 ;
        3445: q <= 32'b00000000000000000000000000000000 ;
        3446: q <= 32'b00000000000000000000000000000000 ;
        3447: q <= 32'b00000000000000000000000000000000 ;
        3448: q <= 32'b00000000000000000000000000000000 ;
        3449: q <= 32'b00000000000000000000000000000000 ;
        3450: q <= 32'b00000000000000000000000000000000 ;
        3451: q <= 32'b00000000000000000000000000000000 ;
        3452: q <= 32'b00000000000000000000000000000000 ;
        3453: q <= 32'b00000000000000000000000000000000 ;
        3454: q <= 32'b00000000000000000000000000000000 ;
        3455: q <= 32'b00000000000000000000000000000000 ;
        3456: q <= 32'b00111100000001110011111110101010 ;
        3457: q <= 32'b10111101101111111000010100000111 ;
        3458: q <= 32'b00111101110100011001000101111011 ;
        3459: q <= 32'b00111101100001100011111111000111 ;
        3460: q <= 32'b10110110001101101011011110001001 ;
        3461: q <= 32'b00111101110011000111010100000010 ;
        3462: q <= 32'b10111101000100111101101011000001 ;
        3463: q <= 32'b00111101001001110010110010101101 ;
        3464: q <= 32'b00111101010010010100100001111101 ;
        3465: q <= 32'b10111101010111000110000000000101 ;
        3466: q <= 32'b10111101101111000101010111000110 ;
        3467: q <= 32'b00111101101011011110000001011001 ;
        3468: q <= 32'b10111101010001011001000000111100 ;
        3469: q <= 32'b00111101101010101110110001011000 ;
        3470: q <= 32'b10111101000111001011000100100110 ;
        3471: q <= 32'b00111011101100001001010110111010 ;
        3472: q <= 32'b00111101000010011001011111101001 ;
        3473: q <= 32'b00111100110101100111110000010110 ;
        3474: q <= 32'b00111101001100101010011110110001 ;
        3475: q <= 32'b00111101010010010011001000101111 ;
        3476: q <= 32'b10111101100001101100010100111000 ;
        3477: q <= 32'b00111101000011000101010010110111 ;
        3478: q <= 32'b00111101101110010111101110110011 ;
        3479: q <= 32'b00111100110100001111101010000011 ;
        3480: q <= 32'b00111101100101001101010101011100 ;
        3481: q <= 32'b10111101101110001001101001111010 ;
        3482: q <= 32'b00111101011111001111100111000010 ;
        3483: q <= 32'b00111101101101100010100110010111 ;
        3484: q <= 32'b00111100110001111101001111011111 ;
        3485: q <= 32'b10111101010100000101101011101000 ;
        3486: q <= 32'b00111010011011110111100111000011 ;
        3487: q <= 32'b00111100100100100000100010100011 ;
        3488: q <= 32'b10111101000111111011100111011000 ;
        3489: q <= 32'b10111100100110101001110011001101 ;
        3490: q <= 32'b00111101010100111111000100110010 ;
        3491: q <= 32'b00111100111111100011111000001110 ;
        3492: q <= 32'b10111101100011001011101011111110 ;
        3493: q <= 32'b10111101011010011011011000011111 ;
        3494: q <= 32'b10111100110011111000110110110111 ;
        3495: q <= 32'b00111011110111000001011000011101 ;
        3496: q <= 32'b10111010110111011111101100011010 ;
        3497: q <= 32'b00111100101101000000001100101001 ;
        3498: q <= 32'b00111101010001000010111111000101 ;
        3499: q <= 32'b10111101011011100010011011111111 ;
        3500: q <= 32'b10111100010110110110111101100001 ;
        3501: q <= 32'b10111100011000110011110100000011 ;
        3502: q <= 32'b10111100111100111000100110000110 ;
        3503: q <= 32'b00111100000111100000000111000101 ;
        3504: q <= 32'b00111101001001001101111010101101 ;
        3505: q <= 32'b00111100110101101000001000110001 ;
        3506: q <= 32'b00111101011111001101110111010000 ;
        3507: q <= 32'b00111100101011001010110111011011 ;
        3508: q <= 32'b00111101100011011100000011010111 ;
        3509: q <= 32'b10111100100101101101100001101100 ;
        3510: q <= 32'b00111100111011000010111000111010 ;
        3511: q <= 32'b10111101101100110011010100100100 ;
        3512: q <= 32'b10111101010110010110100011011010 ;
        3513: q <= 32'b00111101001011110101110101100010 ;
        3514: q <= 32'b00111100010001001010010000100101 ;
        3515: q <= 32'b10111101010100100010001101111011 ;
        3516: q <= 32'b10111100001101100111000101011001 ;
        3517: q <= 32'b00111100110000011110001001101011 ;
        3518: q <= 32'b00111100011010010110011000010010 ;
        3519: q <= 32'b10111101000000001011010101110001 ;
        3520: q <= 32'b10111101000100110011111110011110 ;
        3521: q <= 32'b10111101101100011101101010011000 ;
        3522: q <= 32'b10111101101011101100100000110101 ;
        3523: q <= 32'b10111101101001010010000101110101 ;
        3524: q <= 32'b10111100000111000111110011011110 ;
        3525: q <= 32'b00111101001010011001100000001111 ;
        3526: q <= 32'b10111101001001010000011111010010 ;
        3527: q <= 32'b10111101000110101111110011111000 ;
        3528: q <= 32'b00111101101111000011111011111111 ;
        3529: q <= 32'b00111100110000110010101000010101 ;
        3530: q <= 32'b10111100000111101001000010011110 ;
        3531: q <= 32'b10111101100111001111101101001100 ;
        3532: q <= 32'b00111011100100001010001100010001 ;
        3533: q <= 32'b10111101101111101101111011000011 ;
        3534: q <= 32'b00111101101100000100001110010100 ;
        3535: q <= 32'b00111101101111111110111010010110 ;
        3536: q <= 32'b00111101101100100010110101100100 ;
        3537: q <= 32'b10111101011010001111110000000001 ;
        3538: q <= 32'b10111101110000001000100011001110 ;
        3539: q <= 32'b00111101011100011011001100011110 ;
        3540: q <= 32'b00111101010100010100110010011100 ;
        3541: q <= 32'b10111100101111110111011101010101 ;
        3542: q <= 32'b00111100101000011111001101000000 ;
        3543: q <= 32'b10111101001111010001011110001010 ;
        3544: q <= 32'b00111101100100001111010101010100 ;
        3545: q <= 32'b00111101110010000111001000111100 ;
        3546: q <= 32'b00111101000001010100010111011000 ;
        3547: q <= 32'b10111100101100010011110111111110 ;
        3548: q <= 32'b00111100111101111010100000101101 ;
        3549: q <= 32'b10111100101000110000111001101010 ;
        3550: q <= 32'b00111101100000100011001011010101 ;
        3551: q <= 32'b10111101000010100010111111111001 ;
        3552: q <= 32'b10111101101010001110110000001011 ;
        3553: q <= 32'b00111101001001110101011110010010 ;
        3554: q <= 32'b10111101101100011000011010100111 ;
        3555: q <= 32'b00111100110001010100000010001111 ;
        3556: q <= 32'b00111101101000111101010011010010 ;
        3557: q <= 32'b00111101101010010011010100010011 ;
        3558: q <= 32'b10111101001010101011110010100100 ;
        3559: q <= 32'b10111101011000110011011001111100 ;
        3560: q <= 32'b00000000000000000000000000000000 ;
        3561: q <= 32'b00000000000000000000000000000000 ;
        3562: q <= 32'b00000000000000000000000000000000 ;
        3563: q <= 32'b00000000000000000000000000000000 ;
        3564: q <= 32'b00000000000000000000000000000000 ;
        3565: q <= 32'b00000000000000000000000000000000 ;
        3566: q <= 32'b00000000000000000000000000000000 ;
        3567: q <= 32'b00000000000000000000000000000000 ;
        3568: q <= 32'b00000000000000000000000000000000 ;
        3569: q <= 32'b00000000000000000000000000000000 ;
        3570: q <= 32'b00000000000000000000000000000000 ;
        3571: q <= 32'b00000000000000000000000000000000 ;
        3572: q <= 32'b00000000000000000000000000000000 ;
        3573: q <= 32'b00000000000000000000000000000000 ;
        3574: q <= 32'b00000000000000000000000000000000 ;
        3575: q <= 32'b00000000000000000000000000000000 ;
        3576: q <= 32'b00000000000000000000000000000000 ;
        3577: q <= 32'b00000000000000000000000000000000 ;
        3578: q <= 32'b00000000000000000000000000000000 ;
        3579: q <= 32'b00000000000000000000000000000000 ;
        3580: q <= 32'b00000000000000000000000000000000 ;
        3581: q <= 32'b00000000000000000000000000000000 ;
        3582: q <= 32'b00000000000000000000000000000000 ;
        3583: q <= 32'b00000000000000000000000000000000 ;
        3584: q <= 32'b00111100111000001011101110100101 ;
        3585: q <= 32'b10111100111001011001011010100110 ;
        3586: q <= 32'b00111101100010001010010011111010 ;
        3587: q <= 32'b10111101001110101011010111111001 ;
        3588: q <= 32'b00111101110000100101110110100001 ;
        3589: q <= 32'b00111101100011001000010000100101 ;
        3590: q <= 32'b10111101001000001111100010011111 ;
        3591: q <= 32'b00111101100000000110110110010111 ;
        3592: q <= 32'b00111100010000101110011011001000 ;
        3593: q <= 32'b00111011010000101101000000000100 ;
        3594: q <= 32'b00111101100101011101010100011001 ;
        3595: q <= 32'b10111100111110000000110111010000 ;
        3596: q <= 32'b10111100001001001100000011000011 ;
        3597: q <= 32'b00111101110010001101100010101001 ;
        3598: q <= 32'b00111011010011001101111111000111 ;
        3599: q <= 32'b10111011101110000011001000010100 ;
        3600: q <= 32'b00111101011001100011011101011011 ;
        3601: q <= 32'b00111101001110100110010001010110 ;
        3602: q <= 32'b00111011111000111001101111111010 ;
        3603: q <= 32'b00111011111010010110001011010010 ;
        3604: q <= 32'b10111100110000110011011100010010 ;
        3605: q <= 32'b00111100000111000010111001010111 ;
        3606: q <= 32'b00111101011011101110100100100001 ;
        3607: q <= 32'b00111101010001101011110001111000 ;
        3608: q <= 32'b00111100010100110000101110010110 ;
        3609: q <= 32'b10111101010001000010100000000011 ;
        3610: q <= 32'b00111110000000010111101111110101 ;
        3611: q <= 32'b00111101011001000101111100010110 ;
        3612: q <= 32'b00111101101001101001010101000010 ;
        3613: q <= 32'b10111101101110100001101000010100 ;
        3614: q <= 32'b00111101100000010111110011011101 ;
        3615: q <= 32'b10111101001100110000101111101011 ;
        3616: q <= 32'b00111101011110110100110001011111 ;
        3617: q <= 32'b10111101011011111110001001100011 ;
        3618: q <= 32'b10111101100101001101110111110100 ;
        3619: q <= 32'b00111101011010010110110011100011 ;
        3620: q <= 32'b10111101100100000100011111000101 ;
        3621: q <= 32'b00111101001101001010011100110111 ;
        3622: q <= 32'b00111101011011111000110100000111 ;
        3623: q <= 32'b10111100011010011111011000001100 ;
        3624: q <= 32'b10111101101011000000100001100011 ;
        3625: q <= 32'b10111100101011100101011000000000 ;
        3626: q <= 32'b00111101000011111100011101100101 ;
        3627: q <= 32'b10111101000000010001001110010010 ;
        3628: q <= 32'b00111101110001001011111000010000 ;
        3629: q <= 32'b00111100011100111001010111110110 ;
        3630: q <= 32'b00111100001000110111110101000100 ;
        3631: q <= 32'b00111101100010000010101000010010 ;
        3632: q <= 32'b10111100010001001000000011110101 ;
        3633: q <= 32'b10111100101001011100101000010110 ;
        3634: q <= 32'b00111101011100000010111100001011 ;
        3635: q <= 32'b00111101100010111001101111110010 ;
        3636: q <= 32'b10111101010101011001100010011110 ;
        3637: q <= 32'b10111101011011100111100101011010 ;
        3638: q <= 32'b00111101110001111100110101001110 ;
        3639: q <= 32'b10111101011011110010101001010100 ;
        3640: q <= 32'b00111101101000110010100101101111 ;
        3641: q <= 32'b10111101001111101101010001111010 ;
        3642: q <= 32'b00111011111011000110011100000000 ;
        3643: q <= 32'b00111100101001111111101110001111 ;
        3644: q <= 32'b00111101001101110100111101000101 ;
        3645: q <= 32'b00111101010110001110001100000100 ;
        3646: q <= 32'b10111101000110110110001111101101 ;
        3647: q <= 32'b00111101100001011010000000000100 ;
        3648: q <= 32'b10111101011111100101111100001011 ;
        3649: q <= 32'b00111101011101111010100011011010 ;
        3650: q <= 32'b00111100101111100111100001100110 ;
        3651: q <= 32'b00111101011001110100000111111010 ;
        3652: q <= 32'b10111100110111110000011010101100 ;
        3653: q <= 32'b00111101101101000111101000101011 ;
        3654: q <= 32'b00111101101111010010011011110110 ;
        3655: q <= 32'b00111101101011000101010111011011 ;
        3656: q <= 32'b10111101000111100101101101110111 ;
        3657: q <= 32'b10111101100110101010001110011011 ;
        3658: q <= 32'b00111101110000011010110001001010 ;
        3659: q <= 32'b10111101000100000001111101111101 ;
        3660: q <= 32'b10111011110011001011110001110010 ;
        3661: q <= 32'b00111101011000011100100011101100 ;
        3662: q <= 32'b00111101010110011101001101001100 ;
        3663: q <= 32'b00111101101001100011100000110100 ;
        3664: q <= 32'b00111101000100110100010101001100 ;
        3665: q <= 32'b10111100001110100110011100010100 ;
        3666: q <= 32'b10111101010010001110000101111101 ;
        3667: q <= 32'b00111100011111011001111000110001 ;
        3668: q <= 32'b10111100101001100100110011010111 ;
        3669: q <= 32'b00111101100001101011011101110011 ;
        3670: q <= 32'b10111100000100110001010101100000 ;
        3671: q <= 32'b00111101100000100010101000001010 ;
        3672: q <= 32'b10111101101011010100000100010000 ;
        3673: q <= 32'b10111101001110011101011010110101 ;
        3674: q <= 32'b00111100111101100110011011010100 ;
        3675: q <= 32'b00111101010100101010011000011011 ;
        3676: q <= 32'b10111101110001001111100100101101 ;
        3677: q <= 32'b10111101100000000111011101100010 ;
        3678: q <= 32'b00111101001001010111011000101011 ;
        3679: q <= 32'b00111101010101000110000000000100 ;
        3680: q <= 32'b10111100001100110110110011010101 ;
        3681: q <= 32'b10111101010100110010000000111010 ;
        3682: q <= 32'b00111101001111001000101101101111 ;
        3683: q <= 32'b10111101101010110011010011111100 ;
        3684: q <= 32'b10111101011111011011111101100110 ;
        3685: q <= 32'b10111101011000010110010101110011 ;
        3686: q <= 32'b10111100001010010111010011010101 ;
        3687: q <= 32'b00111100100001111111111001001001 ;
        3688: q <= 32'b00000000000000000000000000000000 ;
        3689: q <= 32'b00000000000000000000000000000000 ;
        3690: q <= 32'b00000000000000000000000000000000 ;
        3691: q <= 32'b00000000000000000000000000000000 ;
        3692: q <= 32'b00000000000000000000000000000000 ;
        3693: q <= 32'b00000000000000000000000000000000 ;
        3694: q <= 32'b00000000000000000000000000000000 ;
        3695: q <= 32'b00000000000000000000000000000000 ;
        3696: q <= 32'b00000000000000000000000000000000 ;
        3697: q <= 32'b00000000000000000000000000000000 ;
        3698: q <= 32'b00000000000000000000000000000000 ;
        3699: q <= 32'b00000000000000000000000000000000 ;
        3700: q <= 32'b00000000000000000000000000000000 ;
        3701: q <= 32'b00000000000000000000000000000000 ;
        3702: q <= 32'b00000000000000000000000000000000 ;
        3703: q <= 32'b00000000000000000000000000000000 ;
        3704: q <= 32'b00000000000000000000000000000000 ;
        3705: q <= 32'b00000000000000000000000000000000 ;
        3706: q <= 32'b00000000000000000000000000000000 ;
        3707: q <= 32'b00000000000000000000000000000000 ;
        3708: q <= 32'b00000000000000000000000000000000 ;
        3709: q <= 32'b00000000000000000000000000000000 ;
        3710: q <= 32'b00000000000000000000000000000000 ;
        3711: q <= 32'b00000000000000000000000000000000 ;
        3712: q <= 32'b10111101110110010110110010101000 ;
        3713: q <= 32'b00111100110101010000011111100011 ;
        3714: q <= 32'b10111101101001110011001101000011 ;
        3715: q <= 32'b10111100001001101101011110100011 ;
        3716: q <= 32'b00111101010010011100001110111100 ;
        3717: q <= 32'b10111101100100000001111100110000 ;
        3718: q <= 32'b10111101010100100011110011111111 ;
        3719: q <= 32'b00111100001010001010000010100011 ;
        3720: q <= 32'b10111101101000101100100100000001 ;
        3721: q <= 32'b10111101100111110101000111100010 ;
        3722: q <= 32'b00111100110010111111110000100001 ;
        3723: q <= 32'b00111101010000000000111001101011 ;
        3724: q <= 32'b00111100111101110011111101011110 ;
        3725: q <= 32'b10111101000001111000001110110000 ;
        3726: q <= 32'b10111101101011011101111110000100 ;
        3727: q <= 32'b10111100110100100101100111011001 ;
        3728: q <= 32'b10111100100000110000011101100101 ;
        3729: q <= 32'b00111101110010011100000110101001 ;
        3730: q <= 32'b00111101010011000010000011001101 ;
        3731: q <= 32'b10111101100001100011000110000101 ;
        3732: q <= 32'b00111101110100010001010100110110 ;
        3733: q <= 32'b10111100001011100001100110100011 ;
        3734: q <= 32'b00111101101100000011101000111010 ;
        3735: q <= 32'b10111101101111000110010010001101 ;
        3736: q <= 32'b00111100101011111111001000111111 ;
        3737: q <= 32'b00111100110011010111000101111001 ;
        3738: q <= 32'b00111011010111110010000100000001 ;
        3739: q <= 32'b10111101001000111100101011110000 ;
        3740: q <= 32'b10111101011000001011011001001000 ;
        3741: q <= 32'b10111101001010010000110001101111 ;
        3742: q <= 32'b10111101001100101010000100010100 ;
        3743: q <= 32'b10111010111001001101111001100111 ;
        3744: q <= 32'b10111101100111010011010011110101 ;
        3745: q <= 32'b00111101010011001010100011111001 ;
        3746: q <= 32'b00111101101110011101010111001010 ;
        3747: q <= 32'b00111100101001111000110001111000 ;
        3748: q <= 32'b00111101101011101010010010110001 ;
        3749: q <= 32'b10111101100001111100110000100111 ;
        3750: q <= 32'b10111101011111000011001111111111 ;
        3751: q <= 32'b00111100111001000110001001101110 ;
        3752: q <= 32'b00111101010101100101000111010101 ;
        3753: q <= 32'b10111100101011111010111011101001 ;
        3754: q <= 32'b00111101101011100100001001110010 ;
        3755: q <= 32'b10111101000110101001101101011101 ;
        3756: q <= 32'b00111101100001111110111101110100 ;
        3757: q <= 32'b10111101100110011111001111001011 ;
        3758: q <= 32'b00111100110100000101001001110000 ;
        3759: q <= 32'b10111101011000000001010001011000 ;
        3760: q <= 32'b10111101000010110101001100100110 ;
        3761: q <= 32'b10111101100110110000111000100001 ;
        3762: q <= 32'b00111100001011001001110001011101 ;
        3763: q <= 32'b10111101110001001001010010101001 ;
        3764: q <= 32'b10111110000010100101010001011111 ;
        3765: q <= 32'b10111100100010011111010001001000 ;
        3766: q <= 32'b00111101001011001010101101000010 ;
        3767: q <= 32'b10111101101111101011010100101001 ;
        3768: q <= 32'b10111101100100011000101010000011 ;
        3769: q <= 32'b00111101100110100011000001110010 ;
        3770: q <= 32'b00111101000100011110110010001000 ;
        3771: q <= 32'b10111101000111111011011101100000 ;
        3772: q <= 32'b00111011100111011111011110000010 ;
        3773: q <= 32'b10111101110011010010011001001000 ;
        3774: q <= 32'b10111101101110110110111000101010 ;
        3775: q <= 32'b10111010011110011001111011100111 ;
        3776: q <= 32'b10111101011001110010010111000001 ;
        3777: q <= 32'b10111101011011010000000010000001 ;
        3778: q <= 32'b10111100101101111010111101001110 ;
        3779: q <= 32'b10111101000000110101011111000110 ;
        3780: q <= 32'b10111101010000100000010010110001 ;
        3781: q <= 32'b00111101001001101101110011000110 ;
        3782: q <= 32'b10111011100001110110100101000011 ;
        3783: q <= 32'b10111101000101101111110000100111 ;
        3784: q <= 32'b10111100001100110011100111111100 ;
        3785: q <= 32'b00111011110000010111110011001110 ;
        3786: q <= 32'b10111101100010000111100100011110 ;
        3787: q <= 32'b10111101011011000000000110000010 ;
        3788: q <= 32'b00111101100010111110101110011010 ;
        3789: q <= 32'b10111101000010001111011101110010 ;
        3790: q <= 32'b00111100100100000011011110101011 ;
        3791: q <= 32'b10111101011011001001111011010001 ;
        3792: q <= 32'b10111101101001001010000010101011 ;
        3793: q <= 32'b00111101100100010101010100000100 ;
        3794: q <= 32'b00111101100011000100011010010111 ;
        3795: q <= 32'b10111101100011000000101101101010 ;
        3796: q <= 32'b00111101100010100111010111101000 ;
        3797: q <= 32'b00111101011101111011011001000001 ;
        3798: q <= 32'b10111101110010000001000111000001 ;
        3799: q <= 32'b10111001111011100111011001010010 ;
        3800: q <= 32'b00111101101010100000011010010010 ;
        3801: q <= 32'b00111101010101111001010101111000 ;
        3802: q <= 32'b10111100001000011100011011011000 ;
        3803: q <= 32'b10111101100111110111000011101011 ;
        3804: q <= 32'b10111101011010101100010011010001 ;
        3805: q <= 32'b00111011010101100110110000100111 ;
        3806: q <= 32'b00111100101011000101100000111001 ;
        3807: q <= 32'b10111101001111101100011011100101 ;
        3808: q <= 32'b10111101100010110100001110100100 ;
        3809: q <= 32'b10111101101101011001010001101001 ;
        3810: q <= 32'b00111101000110000100010101001111 ;
        3811: q <= 32'b10111101100010100011101110001001 ;
        3812: q <= 32'b00111101101100110100010011111110 ;
        3813: q <= 32'b10111101001101011011100100010110 ;
        3814: q <= 32'b10111101011110010100110010101110 ;
        3815: q <= 32'b10111101110000111110111100010010 ;
        3816: q <= 32'b00000000000000000000000000000000 ;
        3817: q <= 32'b00000000000000000000000000000000 ;
        3818: q <= 32'b00000000000000000000000000000000 ;
        3819: q <= 32'b00000000000000000000000000000000 ;
        3820: q <= 32'b00000000000000000000000000000000 ;
        3821: q <= 32'b00000000000000000000000000000000 ;
        3822: q <= 32'b00000000000000000000000000000000 ;
        3823: q <= 32'b00000000000000000000000000000000 ;
        3824: q <= 32'b00000000000000000000000000000000 ;
        3825: q <= 32'b00000000000000000000000000000000 ;
        3826: q <= 32'b00000000000000000000000000000000 ;
        3827: q <= 32'b00000000000000000000000000000000 ;
        3828: q <= 32'b00000000000000000000000000000000 ;
        3829: q <= 32'b00000000000000000000000000000000 ;
        3830: q <= 32'b00000000000000000000000000000000 ;
        3831: q <= 32'b00000000000000000000000000000000 ;
        3832: q <= 32'b00000000000000000000000000000000 ;
        3833: q <= 32'b00000000000000000000000000000000 ;
        3834: q <= 32'b00000000000000000000000000000000 ;
        3835: q <= 32'b00000000000000000000000000000000 ;
        3836: q <= 32'b00000000000000000000000000000000 ;
        3837: q <= 32'b00000000000000000000000000000000 ;
        3838: q <= 32'b00000000000000000000000000000000 ;
        3839: q <= 32'b00000000000000000000000000000000 ;
        3840: q <= 32'b00111101110000011000000100001100 ;
        3841: q <= 32'b00111101110101100110110000110000 ;
        3842: q <= 32'b10111001000001011011111100011100 ;
        3843: q <= 32'b00111101011101100100011001100110 ;
        3844: q <= 32'b00111101101100001110001101000001 ;
        3845: q <= 32'b10111100101001011010100111101011 ;
        3846: q <= 32'b10111011101000110000100010011011 ;
        3847: q <= 32'b00111101011101001010001101000001 ;
        3848: q <= 32'b10111101100011000101101001100000 ;
        3849: q <= 32'b00111100110000000010111011110101 ;
        3850: q <= 32'b00111101110110000011111111111100 ;
        3851: q <= 32'b10111010111000000011001011010100 ;
        3852: q <= 32'b10111101110000101001111110101111 ;
        3853: q <= 32'b10111100111011000001011001010111 ;
        3854: q <= 32'b00111101011010100011011100111100 ;
        3855: q <= 32'b00111101101010110000011011110111 ;
        3856: q <= 32'b00111101000010111111001001101110 ;
        3857: q <= 32'b10111101101000010000110100000111 ;
        3858: q <= 32'b00111100111111000010111100001000 ;
        3859: q <= 32'b00111101111110000110000111001000 ;
        3860: q <= 32'b00111101010110000011001000100000 ;
        3861: q <= 32'b10111100101010110011101111011010 ;
        3862: q <= 32'b10111101011000110100011001111110 ;
        3863: q <= 32'b10111101100110010101011101101111 ;
        3864: q <= 32'b00111101101110100100011111011011 ;
        3865: q <= 32'b00111101011011100100010101101100 ;
        3866: q <= 32'b10111101000011100111010111001100 ;
        3867: q <= 32'b00111110000101100111011011010111 ;
        3868: q <= 32'b00111101110110001100010100000100 ;
        3869: q <= 32'b00111101010010100010111011011110 ;
        3870: q <= 32'b10111101100100001111110100011111 ;
        3871: q <= 32'b10111101010011001010100010110001 ;
        3872: q <= 32'b00111101100111100110001110100000 ;
        3873: q <= 32'b00111101000100111111111111100000 ;
        3874: q <= 32'b10111101110100110010010010011000 ;
        3875: q <= 32'b10111101000111000101001011010011 ;
        3876: q <= 32'b00111101100000111011101110101001 ;
        3877: q <= 32'b10111100101111011110111100111100 ;
        3878: q <= 32'b00111101100101011101110100111101 ;
        3879: q <= 32'b00111101100100110011011000011011 ;
        3880: q <= 32'b10111101110011001011001101010111 ;
        3881: q <= 32'b10111100001100111101000111111001 ;
        3882: q <= 32'b10111101011111110010010101010111 ;
        3883: q <= 32'b00111101001110111110111100010010 ;
        3884: q <= 32'b00111101001001111111010000110111 ;
        3885: q <= 32'b00111110000011011110101101000001 ;
        3886: q <= 32'b10111100100001010010010010100110 ;
        3887: q <= 32'b00111101011110001001111000101010 ;
        3888: q <= 32'b00111101000010111001111011011101 ;
        3889: q <= 32'b10111101010110111011101011111101 ;
        3890: q <= 32'b10111101100010011111101000011010 ;
        3891: q <= 32'b00111101101000011011111011111001 ;
        3892: q <= 32'b00111101101001001100001100000100 ;
        3893: q <= 32'b00111101100010100000000100101000 ;
        3894: q <= 32'b00111100001101111100111100101010 ;
        3895: q <= 32'b10111101001100001011010110110010 ;
        3896: q <= 32'b10111100011101100100101110111100 ;
        3897: q <= 32'b00111100110010100111000000100011 ;
        3898: q <= 32'b10111100100100011101110111100101 ;
        3899: q <= 32'b00111010111000101101010000010011 ;
        3900: q <= 32'b10111101100001110000010000010101 ;
        3901: q <= 32'b00111101111010000100111111001101 ;
        3902: q <= 32'b10111100100101101010101011011010 ;
        3903: q <= 32'b00111101101011111011100111101010 ;
        3904: q <= 32'b00111101001101101001111001000000 ;
        3905: q <= 32'b00111101101001110100110111110011 ;
        3906: q <= 32'b10111101010001000010111011010111 ;
        3907: q <= 32'b10111100001111010010100110001110 ;
        3908: q <= 32'b00111101000001001100100010110000 ;
        3909: q <= 32'b00111101100000101111100100101001 ;
        3910: q <= 32'b10111101000000010100111001000001 ;
        3911: q <= 32'b00111101000101100111111010111100 ;
        3912: q <= 32'b00111101011011101011010010110000 ;
        3913: q <= 32'b00111100101101010100100011001111 ;
        3914: q <= 32'b10111101110001011001011101101010 ;
        3915: q <= 32'b10111101101000101111010110001101 ;
        3916: q <= 32'b10111101011110010101001010101110 ;
        3917: q <= 32'b10111101100111000110010001111111 ;
        3918: q <= 32'b10111101010100000010000000000000 ;
        3919: q <= 32'b00111011111001110010000001000000 ;
        3920: q <= 32'b10111101001110000000100001001000 ;
        3921: q <= 32'b10111101011001010100111010101110 ;
        3922: q <= 32'b10111101010100101100111110111000 ;
        3923: q <= 32'b00111101100010111101000001110100 ;
        3924: q <= 32'b00111101000100000111110010001111 ;
        3925: q <= 32'b10111101101110111101111000001110 ;
        3926: q <= 32'b10111100010000101101000010100100 ;
        3927: q <= 32'b00111101101111011100110001111001 ;
        3928: q <= 32'b00111101110100100100010001111000 ;
        3929: q <= 32'b00111100110110101000110001010001 ;
        3930: q <= 32'b10111001011110100110100110010010 ;
        3931: q <= 32'b10111100000000011000100101010101 ;
        3932: q <= 32'b10111100001100000111100101111111 ;
        3933: q <= 32'b10111101111100001011010101010010 ;
        3934: q <= 32'b00111101100110010010011101110010 ;
        3935: q <= 32'b10111011000011011101110011110010 ;
        3936: q <= 32'b00111101001100111111011000011111 ;
        3937: q <= 32'b00111101101000010011110010010100 ;
        3938: q <= 32'b00111100111110111111111010110001 ;
        3939: q <= 32'b10111100100111011011001100111111 ;
        3940: q <= 32'b10111101100101001001111100101101 ;
        3941: q <= 32'b10111101101000010011111010100011 ;
        3942: q <= 32'b10111100001100100001010101101000 ;
        3943: q <= 32'b10111101100110001101000011000111 ;
        3944: q <= 32'b00000000000000000000000000000000 ;
        3945: q <= 32'b00000000000000000000000000000000 ;
        3946: q <= 32'b00000000000000000000000000000000 ;
        3947: q <= 32'b00000000000000000000000000000000 ;
        3948: q <= 32'b00000000000000000000000000000000 ;
        3949: q <= 32'b00000000000000000000000000000000 ;
        3950: q <= 32'b00000000000000000000000000000000 ;
        3951: q <= 32'b00000000000000000000000000000000 ;
        3952: q <= 32'b00000000000000000000000000000000 ;
        3953: q <= 32'b00000000000000000000000000000000 ;
        3954: q <= 32'b00000000000000000000000000000000 ;
        3955: q <= 32'b00000000000000000000000000000000 ;
        3956: q <= 32'b00000000000000000000000000000000 ;
        3957: q <= 32'b00000000000000000000000000000000 ;
        3958: q <= 32'b00000000000000000000000000000000 ;
        3959: q <= 32'b00000000000000000000000000000000 ;
        3960: q <= 32'b00000000000000000000000000000000 ;
        3961: q <= 32'b00000000000000000000000000000000 ;
        3962: q <= 32'b00000000000000000000000000000000 ;
        3963: q <= 32'b00000000000000000000000000000000 ;
        3964: q <= 32'b00000000000000000000000000000000 ;
        3965: q <= 32'b00000000000000000000000000000000 ;
        3966: q <= 32'b00000000000000000000000000000000 ;
        3967: q <= 32'b00000000000000000000000000000000 ;
        3968: q <= 32'b10111101001111000001100111100000 ;
        3969: q <= 32'b10111101011001001011110110000101 ;
        3970: q <= 32'b10111011111100001111001001100111 ;
        3971: q <= 32'b10111101100000011101101011100011 ;
        3972: q <= 32'b00111101111011001101001100010011 ;
        3973: q <= 32'b00111110000101000111111001111100 ;
        3974: q <= 32'b10111100101111101000001010110000 ;
        3975: q <= 32'b00111101001011101111000111001100 ;
        3976: q <= 32'b10111101010010010011010011001111 ;
        3977: q <= 32'b10111101100111011110011001000111 ;
        3978: q <= 32'b10111011110010000111101101001000 ;
        3979: q <= 32'b00111100101010111011100110100111 ;
        3980: q <= 32'b10111101101011101000110000010111 ;
        3981: q <= 32'b00111101010010010111001101000001 ;
        3982: q <= 32'b10111101010101101110000101110011 ;
        3983: q <= 32'b10111101001010000111100101100001 ;
        3984: q <= 32'b00111110000001001001011011011101 ;
        3985: q <= 32'b00111000100010010011001110110111 ;
        3986: q <= 32'b10111100011111101000001000000110 ;
        3987: q <= 32'b00111011111011101001100001011111 ;
        3988: q <= 32'b10111101000001111010101110101011 ;
        3989: q <= 32'b10111011110111001000010010100111 ;
        3990: q <= 32'b00111101111001100111010100110011 ;
        3991: q <= 32'b10111100000010110010101010001010 ;
        3992: q <= 32'b10111101010000001101101110010110 ;
        3993: q <= 32'b00111101101000110000010000110100 ;
        3994: q <= 32'b00111101100010101111100010111011 ;
        3995: q <= 32'b10111110000110101100101001001100 ;
        3996: q <= 32'b10111101001011000001101100000001 ;
        3997: q <= 32'b10111101101111001101100000011011 ;
        3998: q <= 32'b10111101001001111101011100001100 ;
        3999: q <= 32'b00111100101101111110010101110001 ;
        4000: q <= 32'b00111101001101000111111001011000 ;
        4001: q <= 32'b10111101101010011110010101101011 ;
        4002: q <= 32'b10111100101110001101000000101001 ;
        4003: q <= 32'b10111101101011000001011111111010 ;
        4004: q <= 32'b10111011011011100011110000101011 ;
        4005: q <= 32'b10111101010111001111000000100111 ;
        4006: q <= 32'b00111011010010010011101101001100 ;
        4007: q <= 32'b00111101110100100100111101011110 ;
        4008: q <= 32'b10111101001011010011111111000101 ;
        4009: q <= 32'b10111110000000111110110110110101 ;
        4010: q <= 32'b00111101000001000000110101111101 ;
        4011: q <= 32'b10111101101011011000111100000100 ;
        4012: q <= 32'b00111100101110001100111001100010 ;
        4013: q <= 32'b10111100010110011000111000010001 ;
        4014: q <= 32'b00111011110001011011010001000101 ;
        4015: q <= 32'b00111011011011011100110101001001 ;
        4016: q <= 32'b00111101000000000011101010110111 ;
        4017: q <= 32'b00111100000000101111111110011011 ;
        4018: q <= 32'b00111101100001110111111100010110 ;
        4019: q <= 32'b00111101010101111011100101011101 ;
        4020: q <= 32'b00111101110000000100100111000111 ;
        4021: q <= 32'b00111101100111011010111100101010 ;
        4022: q <= 32'b10111101110010100001110000111110 ;
        4023: q <= 32'b10111101111110000001010100100001 ;
        4024: q <= 32'b00111101110010101000110001000100 ;
        4025: q <= 32'b10111101100000000111110011101000 ;
        4026: q <= 32'b00111101100101110110000111010111 ;
        4027: q <= 32'b00111011001100010100000111100000 ;
        4028: q <= 32'b00111101100001011100100000011100 ;
        4029: q <= 32'b00111101100010101010100001100011 ;
        4030: q <= 32'b10111101101011101110101010111101 ;
        4031: q <= 32'b10111101101000000101011010110010 ;
        4032: q <= 32'b00111101100011001011111100001011 ;
        4033: q <= 32'b00111101010111001110001011101001 ;
        4034: q <= 32'b00111110010100110110010000100000 ;
        4035: q <= 32'b00111101000110111101100111001111 ;
        4036: q <= 32'b00111101010100110101111101011000 ;
        4037: q <= 32'b00111100010111011100011111010001 ;
        4038: q <= 32'b10111100100010001111100101100010 ;
        4039: q <= 32'b10111100100010100001100101111001 ;
        4040: q <= 32'b00111101000010010001111100100011 ;
        4041: q <= 32'b10111101100100010011101000001111 ;
        4042: q <= 32'b00111101111110011100000011001100 ;
        4043: q <= 32'b10111101101001100000000000110001 ;
        4044: q <= 32'b00111101101010111101000100000101 ;
        4045: q <= 32'b10111101100100111000101111100000 ;
        4046: q <= 32'b10111011110100000000111101001010 ;
        4047: q <= 32'b00111110000111111111001010001001 ;
        4048: q <= 32'b10111101011011111010100000010011 ;
        4049: q <= 32'b10111101011001100110101101100011 ;
        4050: q <= 32'b00111100101011000100000011110111 ;
        4051: q <= 32'b10111001001010000110101110100100 ;
        4052: q <= 32'b00111101111001011001000110001110 ;
        4053: q <= 32'b00111101100010101100101011011010 ;
        4054: q <= 32'b10111100101000011101100101011110 ;
        4055: q <= 32'b00111101110010110101111011001000 ;
        4056: q <= 32'b00111101011111100111011111011111 ;
        4057: q <= 32'b10111101000001010111010001111010 ;
        4058: q <= 32'b00111101100000000000001100111110 ;
        4059: q <= 32'b00111101010100101011110010010011 ;
        4060: q <= 32'b00111110011010000101111111011110 ;
        4061: q <= 32'b10111101010010010001111100111110 ;
        4062: q <= 32'b10111101100000001001011100100000 ;
        4063: q <= 32'b10111101001011011110010100100001 ;
        4064: q <= 32'b10111101100011011000110100011111 ;
        4065: q <= 32'b00111101100010001011000101110001 ;
        4066: q <= 32'b00111101001011011001110101001010 ;
        4067: q <= 32'b00111100101110001010110001001011 ;
        4068: q <= 32'b00111101100001000010111110110001 ;
        4069: q <= 32'b10111100111100000100111101110000 ;
        4070: q <= 32'b00111101001000011001110101000000 ;
        4071: q <= 32'b00111101100110100001111010111010 ;
        4072: q <= 32'b00000000000000000000000000000000 ;
        4073: q <= 32'b00000000000000000000000000000000 ;
        4074: q <= 32'b00000000000000000000000000000000 ;
        4075: q <= 32'b00000000000000000000000000000000 ;
        4076: q <= 32'b00000000000000000000000000000000 ;
        4077: q <= 32'b00000000000000000000000000000000 ;
        4078: q <= 32'b00000000000000000000000000000000 ;
        4079: q <= 32'b00000000000000000000000000000000 ;
        4080: q <= 32'b00000000000000000000000000000000 ;
        4081: q <= 32'b00000000000000000000000000000000 ;
        4082: q <= 32'b00000000000000000000000000000000 ;
        4083: q <= 32'b00000000000000000000000000000000 ;
        4084: q <= 32'b00000000000000000000000000000000 ;
        4085: q <= 32'b00000000000000000000000000000000 ;
        4086: q <= 32'b00000000000000000000000000000000 ;
        4087: q <= 32'b00000000000000000000000000000000 ;
        4088: q <= 32'b00000000000000000000000000000000 ;
        4089: q <= 32'b00000000000000000000000000000000 ;
        4090: q <= 32'b00000000000000000000000000000000 ;
        4091: q <= 32'b00000000000000000000000000000000 ;
        4092: q <= 32'b00000000000000000000000000000000 ;
        4093: q <= 32'b00000000000000000000000000000000 ;
        4094: q <= 32'b00000000000000000000000000000000 ;
        4095: q <= 32'b00000000000000000000000000000000 ;
        default: q <= 32'b00000000000000000000000000000000;
    endcase
end

endmodule
