module mem_rom_weight_middle_02 (clock, address, q) ;
parameter DATA_WIDTH =  32;
input clock;
input [11:0] address;
output [DATA_WIDTH-1:0] q;
reg    [DATA_WIDTH-1:0] q;
always@(posedge clock) begin 
    case(address)
        0: q <= 32'b00111100111100000000010111011100 ;
        1: q <= 32'b00111101100111111100101100000110 ;
        2: q <= 32'b10111101011000101110011000001111 ;
        3: q <= 32'b10111101110000001001000000001000 ;
        4: q <= 32'b10111101100011101101000111010000 ;
        5: q <= 32'b00111101000100010011010011001100 ;
        6: q <= 32'b00111100111011100010000101000001 ;
        7: q <= 32'b10111100110111110100000011100000 ;
        8: q <= 32'b00111101011001001011010010000111 ;
        9: q <= 32'b00111101001110111111100001110110 ;
        10: q <= 32'b10111011100110011110000000101011 ;
        11: q <= 32'b00111100000100110011011110110101 ;
        12: q <= 32'b10111101011001010101001000111010 ;
        13: q <= 32'b00111101100011011001110010100111 ;
        14: q <= 32'b10111100110011110111010100101110 ;
        15: q <= 32'b10111100011010000000111111001110 ;
        16: q <= 32'b10111100110011101111111010110110 ;
        17: q <= 32'b00111010011000100111011001111001 ;
        18: q <= 32'b00111101110000011011001001100111 ;
        19: q <= 32'b00111100111111100101000001110011 ;
        20: q <= 32'b10111101010110110001000011001110 ;
        21: q <= 32'b10111101010100000011110000111001 ;
        22: q <= 32'b00111101100011101100000010001010 ;
        23: q <= 32'b10111100111010100010010010111110 ;
        24: q <= 32'b10111100010000001001100001000111 ;
        25: q <= 32'b00111011110001111000110110110101 ;
        26: q <= 32'b00111101010100111110111000011011 ;
        27: q <= 32'b10111100111000010111101001111101 ;
        28: q <= 32'b10111101000101101001111100101010 ;
        29: q <= 32'b10111101101111101110011110111111 ;
        30: q <= 32'b00111101101110101000100111111000 ;
        31: q <= 32'b00111101110100110100110101001110 ;
        32: q <= 32'b00111101110011000011000010001000 ;
        33: q <= 32'b10111101010011000010011011110110 ;
        34: q <= 32'b00111101100111001011111110111110 ;
        35: q <= 32'b10111101010010101100010011101100 ;
        36: q <= 32'b00111101010000001111110011001100 ;
        37: q <= 32'b00111101110011001110001011001110 ;
        38: q <= 32'b10111100101011011001011100011100 ;
        39: q <= 32'b10111101101100111000100001110000 ;
        40: q <= 32'b10111101100010110010000100111010 ;
        41: q <= 32'b00111101100101001100000110010000 ;
        42: q <= 32'b10111101101111111001111010100001 ;
        43: q <= 32'b10111100111101000011111000010011 ;
        44: q <= 32'b10111101000111010000001110111101 ;
        45: q <= 32'b10111011001000100011101111100111 ;
        46: q <= 32'b00111101010011000011101000110100 ;
        47: q <= 32'b00111101100010000001000100000101 ;
        48: q <= 32'b10111100000011010101110111011101 ;
        49: q <= 32'b10111100101101111100011101000110 ;
        50: q <= 32'b00111101000001001110110011010001 ;
        51: q <= 32'b10111101010001000000100010001001 ;
        52: q <= 32'b00111101110011001010000000001111 ;
        53: q <= 32'b10111101011011100011100010101001 ;
        54: q <= 32'b10111101100011101011101011101110 ;
        55: q <= 32'b10111101111000101111100110110011 ;
        56: q <= 32'b00111101100111101111100010101011 ;
        57: q <= 32'b00111110000101110001101110010001 ;
        58: q <= 32'b00111101110100100111010011100001 ;
        59: q <= 32'b10111101001011110000111110110100 ;
        60: q <= 32'b10111101000110110110011110101011 ;
        61: q <= 32'b10111101100111101011111000110011 ;
        62: q <= 32'b10111101101100001100010010101110 ;
        63: q <= 32'b00111101100011011110001001011110 ;
        64: q <= 32'b00111101000110000111100101000010 ;
        65: q <= 32'b10111101001100110101000111100000 ;
        66: q <= 32'b00111100100000000000011110001110 ;
        67: q <= 32'b10111100001010011100110111010010 ;
        68: q <= 32'b00111101101111100110000000000111 ;
        69: q <= 32'b10111101110000001011101010110010 ;
        70: q <= 32'b00111101001100100101010111101000 ;
        71: q <= 32'b00111101100100011010100111111110 ;
        72: q <= 32'b00111100111011111100001110110000 ;
        73: q <= 32'b10111101101101110100001010010100 ;
        74: q <= 32'b10111101000000100100011110100111 ;
        75: q <= 32'b00111101110110010000010110110010 ;
        76: q <= 32'b00111101100110110011000000001011 ;
        77: q <= 32'b00111100110011001000101010110010 ;
        78: q <= 32'b00111101001001110100001110110110 ;
        79: q <= 32'b10111100110000110101101110011001 ;
        80: q <= 32'b00111101000111100000011101110000 ;
        81: q <= 32'b00111101010011011110101111100101 ;
        82: q <= 32'b10111101000001010100011011111001 ;
        83: q <= 32'b00111110000110101110001011100000 ;
        84: q <= 32'b10111101001100100010001101010010 ;
        85: q <= 32'b10111101100111110110111010111010 ;
        86: q <= 32'b00111101100111111110110100010010 ;
        87: q <= 32'b10111101101001101101010011110001 ;
        88: q <= 32'b00111100010101000010110100110100 ;
        89: q <= 32'b10111101100101001010001100001110 ;
        90: q <= 32'b00111101010010000110100001110110 ;
        91: q <= 32'b10111100011100100111001100100000 ;
        92: q <= 32'b10111101100101101011110111101111 ;
        93: q <= 32'b00111101110010110001001010100000 ;
        94: q <= 32'b10111001100100101001011110010010 ;
        95: q <= 32'b10111101010001010001101001100011 ;
        96: q <= 32'b10111101101010100000001111110000 ;
        97: q <= 32'b10111011100000111000001010110011 ;
        98: q <= 32'b00111010000011000001100001011011 ;
        99: q <= 32'b00111100100101010100111101010001 ;
        100: q <= 32'b10111011011110111110010101011111 ;
        101: q <= 32'b00111101100011000010010101000010 ;
        102: q <= 32'b00111101101010100011101100110101 ;
        103: q <= 32'b10111101101011111001100000111100 ;
        104: q <= 32'b00000000000000000000000000000000 ;
        105: q <= 32'b00000000000000000000000000000000 ;
        106: q <= 32'b00000000000000000000000000000000 ;
        107: q <= 32'b00000000000000000000000000000000 ;
        108: q <= 32'b00000000000000000000000000000000 ;
        109: q <= 32'b00000000000000000000000000000000 ;
        110: q <= 32'b00000000000000000000000000000000 ;
        111: q <= 32'b00000000000000000000000000000000 ;
        112: q <= 32'b00000000000000000000000000000000 ;
        113: q <= 32'b00000000000000000000000000000000 ;
        114: q <= 32'b00000000000000000000000000000000 ;
        115: q <= 32'b00000000000000000000000000000000 ;
        116: q <= 32'b00000000000000000000000000000000 ;
        117: q <= 32'b00000000000000000000000000000000 ;
        118: q <= 32'b00000000000000000000000000000000 ;
        119: q <= 32'b00000000000000000000000000000000 ;
        120: q <= 32'b00000000000000000000000000000000 ;
        121: q <= 32'b00000000000000000000000000000000 ;
        122: q <= 32'b00000000000000000000000000000000 ;
        123: q <= 32'b00000000000000000000000000000000 ;
        124: q <= 32'b00000000000000000000000000000000 ;
        125: q <= 32'b00000000000000000000000000000000 ;
        126: q <= 32'b00000000000000000000000000000000 ;
        127: q <= 32'b00000000000000000000000000000000 ;
        128: q <= 32'b00111100001000101110110100100100 ;
        129: q <= 32'b00111110000011011111001001110011 ;
        130: q <= 32'b00111101001000010101010001010010 ;
        131: q <= 32'b10111101100100110001010001100100 ;
        132: q <= 32'b00111100100010100000100110101110 ;
        133: q <= 32'b10111101111110101110010011110011 ;
        134: q <= 32'b10111101100000000101100100101010 ;
        135: q <= 32'b10111101010110000101010110111101 ;
        136: q <= 32'b00111101111001001010001010110011 ;
        137: q <= 32'b00111101100100000001001101010011 ;
        138: q <= 32'b10111110000000110101100100100011 ;
        139: q <= 32'b10111101100001010100010000000001 ;
        140: q <= 32'b10111101101110010001101001010010 ;
        141: q <= 32'b10111100010010101011001000100011 ;
        142: q <= 32'b10111101101010000101011000110010 ;
        143: q <= 32'b00111100101101100110011010100010 ;
        144: q <= 32'b00111101001010000110101111000101 ;
        145: q <= 32'b10111101010001111010111101000010 ;
        146: q <= 32'b10111101011101111100010011100011 ;
        147: q <= 32'b00111101010000010100100010110110 ;
        148: q <= 32'b00111101100100111000101000100110 ;
        149: q <= 32'b10111101001001110110010101100001 ;
        150: q <= 32'b10111100111111011000111110001010 ;
        151: q <= 32'b10111101110011101101010110111010 ;
        152: q <= 32'b00111100111011110100000000111110 ;
        153: q <= 32'b10111101101110100110111111111000 ;
        154: q <= 32'b10111101000111100110000000110100 ;
        155: q <= 32'b10111101000001000010100000111010 ;
        156: q <= 32'b10111101101000000100101000101100 ;
        157: q <= 32'b10111101110000010010010110110001 ;
        158: q <= 32'b00111101101001011000010010101011 ;
        159: q <= 32'b10111100011011100100100000000100 ;
        160: q <= 32'b10111101100101111111010101101011 ;
        161: q <= 32'b00111101000101110001010110110011 ;
        162: q <= 32'b00111101111010001001011001100111 ;
        163: q <= 32'b00111110000000110000000110001111 ;
        164: q <= 32'b00111101001101110011110001100000 ;
        165: q <= 32'b10111101100010101111111110110011 ;
        166: q <= 32'b10111101110010111100101000011101 ;
        167: q <= 32'b10111100101111111111111101001000 ;
        168: q <= 32'b00111101010010101101001111100111 ;
        169: q <= 32'b10111101100011100010100001010011 ;
        170: q <= 32'b00111101000011110000111100101100 ;
        171: q <= 32'b10111010110011100111000011001110 ;
        172: q <= 32'b00111101100111100000010011110100 ;
        173: q <= 32'b00111100111100100101100010011101 ;
        174: q <= 32'b10111101011000010101101011011101 ;
        175: q <= 32'b00111101100011011110110101011111 ;
        176: q <= 32'b10111100101101110001100010110010 ;
        177: q <= 32'b00111101010011111111101010011111 ;
        178: q <= 32'b10111101000111100110101011100010 ;
        179: q <= 32'b10111101011011001110111101000001 ;
        180: q <= 32'b10111101111010101011100100011111 ;
        181: q <= 32'b10111101000110011000010000100000 ;
        182: q <= 32'b10111101001000001111000101011010 ;
        183: q <= 32'b00111100111000110110100000010010 ;
        184: q <= 32'b00111101011101000110101000110000 ;
        185: q <= 32'b10111101101100011001011110101001 ;
        186: q <= 32'b10111101010110011000110110111111 ;
        187: q <= 32'b00111110000000011010010001101010 ;
        188: q <= 32'b00111101101111010000001000010000 ;
        189: q <= 32'b10111101011011101100011100000101 ;
        190: q <= 32'b00111010111010011100011100000100 ;
        191: q <= 32'b00111101010111110011110011110100 ;
        192: q <= 32'b00111010111101011001111001100111 ;
        193: q <= 32'b00111100100001111000000001111100 ;
        194: q <= 32'b10111101101110101101110100110010 ;
        195: q <= 32'b10111100111000110001101101010011 ;
        196: q <= 32'b00111100110000010001010011000010 ;
        197: q <= 32'b10111101001010000010010101000100 ;
        198: q <= 32'b10111101011101001010010110011110 ;
        199: q <= 32'b10111101000000011011100100111110 ;
        200: q <= 32'b00111101100011100100100000001010 ;
        201: q <= 32'b00111101000000110010111001001101 ;
        202: q <= 32'b00111101110000100010100001110100 ;
        203: q <= 32'b00111101011000110110000111000110 ;
        204: q <= 32'b00111101000000011010000011011100 ;
        205: q <= 32'b10111101001111010000101101100100 ;
        206: q <= 32'b00111100001100011011100001111001 ;
        207: q <= 32'b00111101101000110100011111110110 ;
        208: q <= 32'b10111101100110010110100010000011 ;
        209: q <= 32'b00111100000101010001001101011010 ;
        210: q <= 32'b10111101101011001100011010001011 ;
        211: q <= 32'b10111110000000110001000100110111 ;
        212: q <= 32'b10111101011000010100100110111101 ;
        213: q <= 32'b10111101110000011101110011101111 ;
        214: q <= 32'b10111101011111000000010001100010 ;
        215: q <= 32'b10111101100101101101110011010011 ;
        216: q <= 32'b10111101001001110010110110011011 ;
        217: q <= 32'b00111101110001011110100111001010 ;
        218: q <= 32'b00111101101110000011111001110101 ;
        219: q <= 32'b00111101100101010110110001001100 ;
        220: q <= 32'b00111100101111101110011001101100 ;
        221: q <= 32'b00111101110101011110110011000111 ;
        222: q <= 32'b00111110000001001100011001011101 ;
        223: q <= 32'b10111100111001010100001010000101 ;
        224: q <= 32'b00111101010111110011110011010111 ;
        225: q <= 32'b00111101100011000101010111001110 ;
        226: q <= 32'b10111101001001011001111011100000 ;
        227: q <= 32'b00111101010001000111010111010100 ;
        228: q <= 32'b10111100101101100100100100111110 ;
        229: q <= 32'b10111101100000111111101011011100 ;
        230: q <= 32'b10111100010111110111100101111100 ;
        231: q <= 32'b10111101101110111001111001001100 ;
        232: q <= 32'b00000000000000000000000000000000 ;
        233: q <= 32'b00000000000000000000000000000000 ;
        234: q <= 32'b00000000000000000000000000000000 ;
        235: q <= 32'b00000000000000000000000000000000 ;
        236: q <= 32'b00000000000000000000000000000000 ;
        237: q <= 32'b00000000000000000000000000000000 ;
        238: q <= 32'b00000000000000000000000000000000 ;
        239: q <= 32'b00000000000000000000000000000000 ;
        240: q <= 32'b00000000000000000000000000000000 ;
        241: q <= 32'b00000000000000000000000000000000 ;
        242: q <= 32'b00000000000000000000000000000000 ;
        243: q <= 32'b00000000000000000000000000000000 ;
        244: q <= 32'b00000000000000000000000000000000 ;
        245: q <= 32'b00000000000000000000000000000000 ;
        246: q <= 32'b00000000000000000000000000000000 ;
        247: q <= 32'b00000000000000000000000000000000 ;
        248: q <= 32'b00000000000000000000000000000000 ;
        249: q <= 32'b00000000000000000000000000000000 ;
        250: q <= 32'b00000000000000000000000000000000 ;
        251: q <= 32'b00000000000000000000000000000000 ;
        252: q <= 32'b00000000000000000000000000000000 ;
        253: q <= 32'b00000000000000000000000000000000 ;
        254: q <= 32'b00000000000000000000000000000000 ;
        255: q <= 32'b00000000000000000000000000000000 ;
        256: q <= 32'b00111101101100011110001011000010 ;
        257: q <= 32'b00111101100101111011001010110110 ;
        258: q <= 32'b10111101000011001101100000000100 ;
        259: q <= 32'b00111101100100001101000100100010 ;
        260: q <= 32'b00111101111010100110010111101111 ;
        261: q <= 32'b00111101101101011101111110101111 ;
        262: q <= 32'b10111101101100111010011010010001 ;
        263: q <= 32'b00111101110110110100001110100100 ;
        264: q <= 32'b00111100110000111000000011010001 ;
        265: q <= 32'b00111101110101001010010001101110 ;
        266: q <= 32'b10111101010000000101111110001010 ;
        267: q <= 32'b00111100001101100011000011110001 ;
        268: q <= 32'b10111101001110110011101101100011 ;
        269: q <= 32'b10111101000101101011000101001010 ;
        270: q <= 32'b00111011001011010011001001111110 ;
        271: q <= 32'b00111011111101111100110011010111 ;
        272: q <= 32'b10111101101000101000000110101100 ;
        273: q <= 32'b00111101111000010111100111111101 ;
        274: q <= 32'b00111101010011110010100011000110 ;
        275: q <= 32'b10111101010100010101100110101010 ;
        276: q <= 32'b10111011101111111000111110000000 ;
        277: q <= 32'b00111101011100010100101011101000 ;
        278: q <= 32'b10111100110111101111011101101101 ;
        279: q <= 32'b10111101000011010011011110011011 ;
        280: q <= 32'b00111101100100100010000101101011 ;
        281: q <= 32'b00111101000111000101001110010110 ;
        282: q <= 32'b00111100110100010010010011110011 ;
        283: q <= 32'b00111100000010101000100000100111 ;
        284: q <= 32'b10111101100100000110010010110001 ;
        285: q <= 32'b10111101000110100011101000010110 ;
        286: q <= 32'b00111110000010111011011101000101 ;
        287: q <= 32'b00111100100111111000110010101111 ;
        288: q <= 32'b00111100011110010100011000001111 ;
        289: q <= 32'b00111100010001011111110011001011 ;
        290: q <= 32'b10111101101011110110011010000011 ;
        291: q <= 32'b00111101001101111110100101011011 ;
        292: q <= 32'b10111101010111011000011111101111 ;
        293: q <= 32'b00111100011011101011000000000010 ;
        294: q <= 32'b00111101010110001011110000100100 ;
        295: q <= 32'b10111101010110100011000010110101 ;
        296: q <= 32'b00111011101011100101010111001110 ;
        297: q <= 32'b10111100111101001110001010101010 ;
        298: q <= 32'b10111101101000100100001000011011 ;
        299: q <= 32'b00111101101100110110001110100000 ;
        300: q <= 32'b10111100110110111111111010110100 ;
        301: q <= 32'b10111101101011110011111100001010 ;
        302: q <= 32'b00111101011111111100010000010000 ;
        303: q <= 32'b00111101001011000100001011011011 ;
        304: q <= 32'b10111110000011000001010001110000 ;
        305: q <= 32'b10111011111000001100111100100100 ;
        306: q <= 32'b00111100010111001011110011101110 ;
        307: q <= 32'b10111101001011010000001001000001 ;
        308: q <= 32'b10111101100110000111100101000110 ;
        309: q <= 32'b00111101111011110101111010101101 ;
        310: q <= 32'b10111101110101100010111110101001 ;
        311: q <= 32'b00111101000000000011010010011100 ;
        312: q <= 32'b00111110000111011111101000010001 ;
        313: q <= 32'b00111101101101001000101111100000 ;
        314: q <= 32'b10111101001101100101101110011011 ;
        315: q <= 32'b00111101110000101101110010111000 ;
        316: q <= 32'b00111101011100001001011010100100 ;
        317: q <= 32'b10111100100100110010100001001010 ;
        318: q <= 32'b00111101000100010101101011011111 ;
        319: q <= 32'b00111101101000010100001000011110 ;
        320: q <= 32'b00111101000011000001000011100001 ;
        321: q <= 32'b00111101010111001101111100101010 ;
        322: q <= 32'b00111101000011000101111000000111 ;
        323: q <= 32'b10111100110111001110110111000111 ;
        324: q <= 32'b00111101011110000000011100010110 ;
        325: q <= 32'b10111101011111111110001010110011 ;
        326: q <= 32'b10111101101111010010101000101110 ;
        327: q <= 32'b10111101000001011111010010100110 ;
        328: q <= 32'b00111100101110100001111111000000 ;
        329: q <= 32'b10111100011110001110001110000010 ;
        330: q <= 32'b00111101100100100101111000101000 ;
        331: q <= 32'b10111101110000001000001010011110 ;
        332: q <= 32'b10111100000011111101001000100101 ;
        333: q <= 32'b00111101100110110111001000111100 ;
        334: q <= 32'b00111101101000111000010101110100 ;
        335: q <= 32'b00111101001111011111111101101110 ;
        336: q <= 32'b10111110000110100000010111110000 ;
        337: q <= 32'b00111100111101100011110111101001 ;
        338: q <= 32'b00111101110000001110011100111010 ;
        339: q <= 32'b10111101101001000111110100001000 ;
        340: q <= 32'b00111110000000001001001110110011 ;
        341: q <= 32'b00111101011001001000000001001001 ;
        342: q <= 32'b10111101101000011011001110000111 ;
        343: q <= 32'b00111100101110010100100010101110 ;
        344: q <= 32'b00111101011111110011001011101010 ;
        345: q <= 32'b00111101010110100000101011011110 ;
        346: q <= 32'b10111101000000010100111010111011 ;
        347: q <= 32'b10111101001010101101101101101101 ;
        348: q <= 32'b10111100111000010000011000001000 ;
        349: q <= 32'b10111101000110101101100000111000 ;
        350: q <= 32'b00111100100010110111000100111011 ;
        351: q <= 32'b10111100001011111110110010000101 ;
        352: q <= 32'b10111101100100010011110001100111 ;
        353: q <= 32'b00111101011000010100010101011010 ;
        354: q <= 32'b10111100100000000000001101110111 ;
        355: q <= 32'b00111101000011100101010101101010 ;
        356: q <= 32'b10111101110100011010100101010111 ;
        357: q <= 32'b10111011101110001010010101101110 ;
        358: q <= 32'b10111100101110100000001001010111 ;
        359: q <= 32'b10111101101011101010011101000001 ;
        360: q <= 32'b00000000000000000000000000000000 ;
        361: q <= 32'b00000000000000000000000000000000 ;
        362: q <= 32'b00000000000000000000000000000000 ;
        363: q <= 32'b00000000000000000000000000000000 ;
        364: q <= 32'b00000000000000000000000000000000 ;
        365: q <= 32'b00000000000000000000000000000000 ;
        366: q <= 32'b00000000000000000000000000000000 ;
        367: q <= 32'b00000000000000000000000000000000 ;
        368: q <= 32'b00000000000000000000000000000000 ;
        369: q <= 32'b00000000000000000000000000000000 ;
        370: q <= 32'b00000000000000000000000000000000 ;
        371: q <= 32'b00000000000000000000000000000000 ;
        372: q <= 32'b00000000000000000000000000000000 ;
        373: q <= 32'b00000000000000000000000000000000 ;
        374: q <= 32'b00000000000000000000000000000000 ;
        375: q <= 32'b00000000000000000000000000000000 ;
        376: q <= 32'b00000000000000000000000000000000 ;
        377: q <= 32'b00000000000000000000000000000000 ;
        378: q <= 32'b00000000000000000000000000000000 ;
        379: q <= 32'b00000000000000000000000000000000 ;
        380: q <= 32'b00000000000000000000000000000000 ;
        381: q <= 32'b00000000000000000000000000000000 ;
        382: q <= 32'b00000000000000000000000000000000 ;
        383: q <= 32'b00000000000000000000000000000000 ;
        384: q <= 32'b00111101100011000100101000010000 ;
        385: q <= 32'b10111100100000001100111101100111 ;
        386: q <= 32'b10111101011111001101100001001000 ;
        387: q <= 32'b00111110000001001001000011011100 ;
        388: q <= 32'b10111101000010011100011111110000 ;
        389: q <= 32'b10111101000110110001111011000101 ;
        390: q <= 32'b00111101110001001010010111111010 ;
        391: q <= 32'b00111101101001100101110100110001 ;
        392: q <= 32'b10111101010100000001001000011011 ;
        393: q <= 32'b00111101110101011001110101111101 ;
        394: q <= 32'b10111011111111001000100001000010 ;
        395: q <= 32'b10111101011111001100101110010111 ;
        396: q <= 32'b00111010100000110010000011010010 ;
        397: q <= 32'b10111100100111011011110110101000 ;
        398: q <= 32'b10111101010000010111110110111111 ;
        399: q <= 32'b00111100100010001011000011101100 ;
        400: q <= 32'b10111101101000010010100001101111 ;
        401: q <= 32'b00111100101110111110000110010110 ;
        402: q <= 32'b00111101001100100001100000101001 ;
        403: q <= 32'b00111100011111001110000101011101 ;
        404: q <= 32'b10111101111000010001101000000001 ;
        405: q <= 32'b10111101001111110011010110010001 ;
        406: q <= 32'b10111101010000000001111001001010 ;
        407: q <= 32'b10111101000101011101010001101001 ;
        408: q <= 32'b00111101100011110001011001100100 ;
        409: q <= 32'b00111100001101011000000111001000 ;
        410: q <= 32'b00111101000101011010010001100110 ;
        411: q <= 32'b00111101011101101000101100101111 ;
        412: q <= 32'b10111101101110010010001010011111 ;
        413: q <= 32'b10111101000111100000111110110011 ;
        414: q <= 32'b00111101101101011111101111000010 ;
        415: q <= 32'b00111101100110001000000111101101 ;
        416: q <= 32'b00111101000000110110001110000100 ;
        417: q <= 32'b10111101000000010001110001000001 ;
        418: q <= 32'b10111101101111101001001011110100 ;
        419: q <= 32'b10111101011001110101010100111101 ;
        420: q <= 32'b10111100100110010110000010110001 ;
        421: q <= 32'b00111101010101001101011110001101 ;
        422: q <= 32'b10111100101010110010111010001010 ;
        423: q <= 32'b10111101111000111011011110101110 ;
        424: q <= 32'b10111011101000000100110011001101 ;
        425: q <= 32'b10111101110100111100011001011000 ;
        426: q <= 32'b10111101100100111001110111101110 ;
        427: q <= 32'b00111101100110101010100001110111 ;
        428: q <= 32'b00111101101011011100111110100101 ;
        429: q <= 32'b00111101101101111011011110100111 ;
        430: q <= 32'b10111100111110110100110110101101 ;
        431: q <= 32'b00111101111010110111011101111110 ;
        432: q <= 32'b10111101101000000011101100110101 ;
        433: q <= 32'b00111101101010100110110000110001 ;
        434: q <= 32'b00111100111111110100111011011000 ;
        435: q <= 32'b00111101110000100011011010101100 ;
        436: q <= 32'b10111101010011001111011010111001 ;
        437: q <= 32'b10111101100101001000000010111001 ;
        438: q <= 32'b10111101111011101111110001011101 ;
        439: q <= 32'b00111101010111010111001110101000 ;
        440: q <= 32'b10111100110101101011001010001101 ;
        441: q <= 32'b00111101011111010100100010110010 ;
        442: q <= 32'b00111101100011100110111110101000 ;
        443: q <= 32'b10111101100000010011010101111110 ;
        444: q <= 32'b10111011010011001111110100001010 ;
        445: q <= 32'b00111100111100110010011110001001 ;
        446: q <= 32'b00111101100011100001100111010100 ;
        447: q <= 32'b10111100101010011001011011110010 ;
        448: q <= 32'b10111100101110010010001011111000 ;
        449: q <= 32'b00111011110111101000011101011101 ;
        450: q <= 32'b00111100011000010101001110000011 ;
        451: q <= 32'b10111101001000001110110010111011 ;
        452: q <= 32'b00111101010011111110110110101101 ;
        453: q <= 32'b00111101001011011011100011000110 ;
        454: q <= 32'b10111011100011100100111110111011 ;
        455: q <= 32'b00111101101011110110001111011011 ;
        456: q <= 32'b00111100101111100010000100110100 ;
        457: q <= 32'b00111101101001111111100001000111 ;
        458: q <= 32'b00111101100101011000010101011100 ;
        459: q <= 32'b10111101110100000010100100101100 ;
        460: q <= 32'b10111101100011010000111001001000 ;
        461: q <= 32'b10111101000101001110001110100001 ;
        462: q <= 32'b00111101010111100110011010111011 ;
        463: q <= 32'b10111100001000100000000011110000 ;
        464: q <= 32'b10111100111001000000110011011101 ;
        465: q <= 32'b00111110000001000111011001001000 ;
        466: q <= 32'b10111100101110001100011010000001 ;
        467: q <= 32'b00111101100000111100110000010111 ;
        468: q <= 32'b00111101100010100111101001101101 ;
        469: q <= 32'b00111101100001001110011001001101 ;
        470: q <= 32'b00111001011101010110010000101001 ;
        471: q <= 32'b00111100010010110101001010001001 ;
        472: q <= 32'b10111101001011010011111001101110 ;
        473: q <= 32'b00111101011100111000111011111000 ;
        474: q <= 32'b00111101101101111011000111111010 ;
        475: q <= 32'b10111101100100111001111101101100 ;
        476: q <= 32'b00111101010010010101110000100101 ;
        477: q <= 32'b00111010111001011010011011010111 ;
        478: q <= 32'b00111011100001110110110011101101 ;
        479: q <= 32'b00111100100000001011111100101010 ;
        480: q <= 32'b10111101101010000010001011000110 ;
        481: q <= 32'b10111100111111111101001101000111 ;
        482: q <= 32'b00111100000110111101100001111111 ;
        483: q <= 32'b10111101011000101001011000100101 ;
        484: q <= 32'b00111101011001100111111000110000 ;
        485: q <= 32'b10111101101011100000000001001011 ;
        486: q <= 32'b00111100000100100001100010011111 ;
        487: q <= 32'b00111101000011100110010011110011 ;
        488: q <= 32'b00000000000000000000000000000000 ;
        489: q <= 32'b00000000000000000000000000000000 ;
        490: q <= 32'b00000000000000000000000000000000 ;
        491: q <= 32'b00000000000000000000000000000000 ;
        492: q <= 32'b00000000000000000000000000000000 ;
        493: q <= 32'b00000000000000000000000000000000 ;
        494: q <= 32'b00000000000000000000000000000000 ;
        495: q <= 32'b00000000000000000000000000000000 ;
        496: q <= 32'b00000000000000000000000000000000 ;
        497: q <= 32'b00000000000000000000000000000000 ;
        498: q <= 32'b00000000000000000000000000000000 ;
        499: q <= 32'b00000000000000000000000000000000 ;
        500: q <= 32'b00000000000000000000000000000000 ;
        501: q <= 32'b00000000000000000000000000000000 ;
        502: q <= 32'b00000000000000000000000000000000 ;
        503: q <= 32'b00000000000000000000000000000000 ;
        504: q <= 32'b00000000000000000000000000000000 ;
        505: q <= 32'b00000000000000000000000000000000 ;
        506: q <= 32'b00000000000000000000000000000000 ;
        507: q <= 32'b00000000000000000000000000000000 ;
        508: q <= 32'b00000000000000000000000000000000 ;
        509: q <= 32'b00000000000000000000000000000000 ;
        510: q <= 32'b00000000000000000000000000000000 ;
        511: q <= 32'b00000000000000000000000000000000 ;
        512: q <= 32'b00111101111000010101101000011001 ;
        513: q <= 32'b00111101100110110000000101111000 ;
        514: q <= 32'b00111101101000110001011110010100 ;
        515: q <= 32'b00111100101011011010101011110011 ;
        516: q <= 32'b00111101101101001101001001011010 ;
        517: q <= 32'b00111101000000001011010100010011 ;
        518: q <= 32'b10111101001100010000100111101011 ;
        519: q <= 32'b10111101100011110010000111110111 ;
        520: q <= 32'b00111101010011101001110111111010 ;
        521: q <= 32'b10111100111110001011000000101100 ;
        522: q <= 32'b10111101101000001000101110111001 ;
        523: q <= 32'b00111100001000110101011010000001 ;
        524: q <= 32'b00111101011111101010111010111100 ;
        525: q <= 32'b10111101011000101010111100010011 ;
        526: q <= 32'b00111101011010011100011111111001 ;
        527: q <= 32'b10111101000001110101010010010011 ;
        528: q <= 32'b10111100111101001101001011011111 ;
        529: q <= 32'b10111101110010011000011100011000 ;
        530: q <= 32'b10111101100100110010110011110001 ;
        531: q <= 32'b10111101010011001110111110001100 ;
        532: q <= 32'b10111101001000011011010111000110 ;
        533: q <= 32'b00111100010110111100000000101010 ;
        534: q <= 32'b00111101101011100100101000100011 ;
        535: q <= 32'b00111010111100111000011010010001 ;
        536: q <= 32'b10111100101000001100100011101111 ;
        537: q <= 32'b10111101001000100101001110001111 ;
        538: q <= 32'b00111101010000000101100001000001 ;
        539: q <= 32'b10111000100000010001110110100001 ;
        540: q <= 32'b10111100110100010100100011110100 ;
        541: q <= 32'b10111101001100110001111011001111 ;
        542: q <= 32'b10111100110111010110111010011011 ;
        543: q <= 32'b00111101000100111001100010010101 ;
        544: q <= 32'b00111101010100111011111000110100 ;
        545: q <= 32'b00111100110101100001000000000011 ;
        546: q <= 32'b00111101000001110000000110111111 ;
        547: q <= 32'b00111100110100101101010000110110 ;
        548: q <= 32'b10111101100110010000011010111000 ;
        549: q <= 32'b00111101100101001011111111010000 ;
        550: q <= 32'b00111100101110101010011101100000 ;
        551: q <= 32'b00111101001010100110011100111011 ;
        552: q <= 32'b10111101000010101000010101000110 ;
        553: q <= 32'b00111101001010001100001111100000 ;
        554: q <= 32'b10111100110101000110011111011001 ;
        555: q <= 32'b00111101010111000010100100010111 ;
        556: q <= 32'b00111101011001100000000001010100 ;
        557: q <= 32'b10111011100100011011000110011110 ;
        558: q <= 32'b00111011100001110111001100001011 ;
        559: q <= 32'b10111100111000000110001101111011 ;
        560: q <= 32'b10111101000111010110011111000110 ;
        561: q <= 32'b10111100111010010111101001001111 ;
        562: q <= 32'b10111101011111110011101000101100 ;
        563: q <= 32'b10111101101110010111000001011110 ;
        564: q <= 32'b00111101111101111100110001101111 ;
        565: q <= 32'b00111101100101011111111000010101 ;
        566: q <= 32'b00111101111010001010101000100100 ;
        567: q <= 32'b00111101101010010101011101001110 ;
        568: q <= 32'b00111101100000000011000011101101 ;
        569: q <= 32'b00111101110001010110101001011010 ;
        570: q <= 32'b00111101001100011010000010011001 ;
        571: q <= 32'b00111101100001111111100001001100 ;
        572: q <= 32'b00111100111010110000110111010101 ;
        573: q <= 32'b00111101000110011101110001101111 ;
        574: q <= 32'b00111011011100010101101110111111 ;
        575: q <= 32'b00111101000111010100000010101000 ;
        576: q <= 32'b10111100100111100011100011111011 ;
        577: q <= 32'b00111101000101100000111111100001 ;
        578: q <= 32'b00111100001011111011110100010011 ;
        579: q <= 32'b00111101010100000110111111110000 ;
        580: q <= 32'b10111101100011001000010000011111 ;
        581: q <= 32'b00111011011000111111000010100110 ;
        582: q <= 32'b10111101011110000001010001111101 ;
        583: q <= 32'b00111100010000100111110010111010 ;
        584: q <= 32'b00111100000110010110011111010111 ;
        585: q <= 32'b10111101010101100111011111010000 ;
        586: q <= 32'b10111101100011111000000010000111 ;
        587: q <= 32'b00111101100100100100100100100100 ;
        588: q <= 32'b00111101010111111100110011110011 ;
        589: q <= 32'b00111101001011111101110001001111 ;
        590: q <= 32'b00111100011101100101111001001101 ;
        591: q <= 32'b10111101000101001100111011101100 ;
        592: q <= 32'b00111101011101111010010000111101 ;
        593: q <= 32'b10111101100111111010001110100111 ;
        594: q <= 32'b00111100011101011001011100111111 ;
        595: q <= 32'b10111101001000011101001100111101 ;
        596: q <= 32'b00111101000110010100110111011000 ;
        597: q <= 32'b10111100101101010110010100010000 ;
        598: q <= 32'b00111101100100011000101001010101 ;
        599: q <= 32'b10111101100111010000011000011001 ;
        600: q <= 32'b00111101101011100100000001001110 ;
        601: q <= 32'b00111101110001101010101101011011 ;
        602: q <= 32'b00111011110100110001111110010001 ;
        603: q <= 32'b00111011100011001001110010100110 ;
        604: q <= 32'b10111101110010100101100001000010 ;
        605: q <= 32'b00111011001000001101100001110011 ;
        606: q <= 32'b10111101100001011011011011000101 ;
        607: q <= 32'b10111101100110011111011111010111 ;
        608: q <= 32'b10111100011000011100100100101001 ;
        609: q <= 32'b00111101110000011101001000111010 ;
        610: q <= 32'b10111011010001100000001101111001 ;
        611: q <= 32'b10111101001010001100110011011000 ;
        612: q <= 32'b10111101000000100011100011110100 ;
        613: q <= 32'b00111101101110011000011111011111 ;
        614: q <= 32'b10111101101101100100100110000111 ;
        615: q <= 32'b10111101100110001100110101100010 ;
        616: q <= 32'b00000000000000000000000000000000 ;
        617: q <= 32'b00000000000000000000000000000000 ;
        618: q <= 32'b00000000000000000000000000000000 ;
        619: q <= 32'b00000000000000000000000000000000 ;
        620: q <= 32'b00000000000000000000000000000000 ;
        621: q <= 32'b00000000000000000000000000000000 ;
        622: q <= 32'b00000000000000000000000000000000 ;
        623: q <= 32'b00000000000000000000000000000000 ;
        624: q <= 32'b00000000000000000000000000000000 ;
        625: q <= 32'b00000000000000000000000000000000 ;
        626: q <= 32'b00000000000000000000000000000000 ;
        627: q <= 32'b00000000000000000000000000000000 ;
        628: q <= 32'b00000000000000000000000000000000 ;
        629: q <= 32'b00000000000000000000000000000000 ;
        630: q <= 32'b00000000000000000000000000000000 ;
        631: q <= 32'b00000000000000000000000000000000 ;
        632: q <= 32'b00000000000000000000000000000000 ;
        633: q <= 32'b00000000000000000000000000000000 ;
        634: q <= 32'b00000000000000000000000000000000 ;
        635: q <= 32'b00000000000000000000000000000000 ;
        636: q <= 32'b00000000000000000000000000000000 ;
        637: q <= 32'b00000000000000000000000000000000 ;
        638: q <= 32'b00000000000000000000000000000000 ;
        639: q <= 32'b00000000000000000000000000000000 ;
        640: q <= 32'b00111101110001100110000011101000 ;
        641: q <= 32'b00111011100010101111001101111110 ;
        642: q <= 32'b00111110001001101011010000110010 ;
        643: q <= 32'b10111101000001010011100000111001 ;
        644: q <= 32'b10111101101110010100001010100110 ;
        645: q <= 32'b00111101011100011110101101001101 ;
        646: q <= 32'b00111101100000110101110111111101 ;
        647: q <= 32'b00111101011110110111010011100010 ;
        648: q <= 32'b10111101110001111110011110001010 ;
        649: q <= 32'b10111100010001111100011010110000 ;
        650: q <= 32'b10111101101111011110111100011101 ;
        651: q <= 32'b10111011111001100110101100000110 ;
        652: q <= 32'b00111101101011110011010111011101 ;
        653: q <= 32'b00111100100010101010010011101010 ;
        654: q <= 32'b00111110000010111101000100110100 ;
        655: q <= 32'b10111101011111110110000001010111 ;
        656: q <= 32'b10111110000101000000111010111001 ;
        657: q <= 32'b10111101100001010011010111010000 ;
        658: q <= 32'b00111110001010001100110001011110 ;
        659: q <= 32'b00111101001101101001001101101100 ;
        660: q <= 32'b00111100001101011000100000110000 ;
        661: q <= 32'b00111100101111011111010101010110 ;
        662: q <= 32'b10111100101111101011100110001011 ;
        663: q <= 32'b00111110001001010011001001000111 ;
        664: q <= 32'b00111101101011101011000111010101 ;
        665: q <= 32'b10111100100110011110101010101111 ;
        666: q <= 32'b10111011110101001011000100100001 ;
        667: q <= 32'b10111101011011110100000100100111 ;
        668: q <= 32'b00111110000011001101001101001101 ;
        669: q <= 32'b10111101101100010100010101101100 ;
        670: q <= 32'b10111101111010111011110111011101 ;
        671: q <= 32'b00111101101111101000100011100011 ;
        672: q <= 32'b00111100111001011110111101100011 ;
        673: q <= 32'b00111101011000011000110000100001 ;
        674: q <= 32'b00111101001010010100111001010001 ;
        675: q <= 32'b10111100011011101011110011111101 ;
        676: q <= 32'b00111101011010010010010111000110 ;
        677: q <= 32'b10111101000001011100110101010111 ;
        678: q <= 32'b00111101011010010001111111000111 ;
        679: q <= 32'b00111110000110010100110011101001 ;
        680: q <= 32'b10111100101100110101011111110100 ;
        681: q <= 32'b00111011110110000111010011101100 ;
        682: q <= 32'b00111101100111101101111111011010 ;
        683: q <= 32'b10111110001001101010010111010111 ;
        684: q <= 32'b10111100110001010000101010011110 ;
        685: q <= 32'b00111101010011111011011000010001 ;
        686: q <= 32'b10111101100100110101011110111001 ;
        687: q <= 32'b00111101000101100001001011110110 ;
        688: q <= 32'b00111011011000001001101010101001 ;
        689: q <= 32'b00111101001101100100011000101010 ;
        690: q <= 32'b10111101100110111000000000110111 ;
        691: q <= 32'b00111101011110111111111111111010 ;
        692: q <= 32'b10111101010000110100111010100010 ;
        693: q <= 32'b00111101010110110010111101011111 ;
        694: q <= 32'b00111101101000000101010100011100 ;
        695: q <= 32'b00111100110100101111010000010010 ;
        696: q <= 32'b00111101001111101010001101101011 ;
        697: q <= 32'b00111101001000111001001110001101 ;
        698: q <= 32'b10111101000000110011100101100100 ;
        699: q <= 32'b10111101101001001000100010011111 ;
        700: q <= 32'b00111101110001000111011010001000 ;
        701: q <= 32'b10111101010100111001101110011010 ;
        702: q <= 32'b10111101011011001010011101010110 ;
        703: q <= 32'b10111100100110001100101011100001 ;
        704: q <= 32'b00111101000001000011010100000101 ;
        705: q <= 32'b00111100011001010111101101110011 ;
        706: q <= 32'b10111010011001111110011010010011 ;
        707: q <= 32'b10111100000001110111000001111101 ;
        708: q <= 32'b00111101101110001101001010110011 ;
        709: q <= 32'b00111101110010011000101110110110 ;
        710: q <= 32'b00111101100011010100000100011011 ;
        711: q <= 32'b10111101110111111111000100100010 ;
        712: q <= 32'b00111101000010101011000110100000 ;
        713: q <= 32'b10111101001010001101110110100000 ;
        714: q <= 32'b00111101100011011110010111110110 ;
        715: q <= 32'b10111101010100000100000001001000 ;
        716: q <= 32'b00111100001110001011110010100101 ;
        717: q <= 32'b00111101010000100000000100000101 ;
        718: q <= 32'b10111100011010110001011011101000 ;
        719: q <= 32'b00111110011010100010100100111010 ;
        720: q <= 32'b10111101011010011001101010001010 ;
        721: q <= 32'b10111101111000111001111011011100 ;
        722: q <= 32'b10111100101010110101111101111000 ;
        723: q <= 32'b00111101111000100010000010000110 ;
        724: q <= 32'b00111100100011001111000010100001 ;
        725: q <= 32'b10111101110011110000100111011010 ;
        726: q <= 32'b00111100100010110010101000010110 ;
        727: q <= 32'b00111101100110101001110000010110 ;
        728: q <= 32'b00111100100000000000101001101111 ;
        729: q <= 32'b10111101000011110101110111011010 ;
        730: q <= 32'b00111101010010000011011010011010 ;
        731: q <= 32'b00111101110001111111100000011010 ;
        732: q <= 32'b00111101110010010110110101111101 ;
        733: q <= 32'b10111101011110101010011011011110 ;
        734: q <= 32'b10111101000000111001001011011101 ;
        735: q <= 32'b00111100110101100111100001100100 ;
        736: q <= 32'b10111010101001001111011010000101 ;
        737: q <= 32'b00111101100000101011111011000111 ;
        738: q <= 32'b10111101010011001110000101011110 ;
        739: q <= 32'b00111100111000101111111001101101 ;
        740: q <= 32'b00111101011001111101001001110000 ;
        741: q <= 32'b10111101011111101001110010101100 ;
        742: q <= 32'b00111101101110110010110011111000 ;
        743: q <= 32'b00111101101001000000001111010111 ;
        744: q <= 32'b00000000000000000000000000000000 ;
        745: q <= 32'b00000000000000000000000000000000 ;
        746: q <= 32'b00000000000000000000000000000000 ;
        747: q <= 32'b00000000000000000000000000000000 ;
        748: q <= 32'b00000000000000000000000000000000 ;
        749: q <= 32'b00000000000000000000000000000000 ;
        750: q <= 32'b00000000000000000000000000000000 ;
        751: q <= 32'b00000000000000000000000000000000 ;
        752: q <= 32'b00000000000000000000000000000000 ;
        753: q <= 32'b00000000000000000000000000000000 ;
        754: q <= 32'b00000000000000000000000000000000 ;
        755: q <= 32'b00000000000000000000000000000000 ;
        756: q <= 32'b00000000000000000000000000000000 ;
        757: q <= 32'b00000000000000000000000000000000 ;
        758: q <= 32'b00000000000000000000000000000000 ;
        759: q <= 32'b00000000000000000000000000000000 ;
        760: q <= 32'b00000000000000000000000000000000 ;
        761: q <= 32'b00000000000000000000000000000000 ;
        762: q <= 32'b00000000000000000000000000000000 ;
        763: q <= 32'b00000000000000000000000000000000 ;
        764: q <= 32'b00000000000000000000000000000000 ;
        765: q <= 32'b00000000000000000000000000000000 ;
        766: q <= 32'b00000000000000000000000000000000 ;
        767: q <= 32'b00000000000000000000000000000000 ;
        768: q <= 32'b10111101001100110010100111001110 ;
        769: q <= 32'b00111011110001011111111001100100 ;
        770: q <= 32'b10111101000010011010010100111011 ;
        771: q <= 32'b10111101001100011010101100100101 ;
        772: q <= 32'b00111100001110011000010110110010 ;
        773: q <= 32'b00111100100011001100001111010010 ;
        774: q <= 32'b10111101110100111000110010100000 ;
        775: q <= 32'b10111101001101110101111000101110 ;
        776: q <= 32'b00111101110000110010110001011110 ;
        777: q <= 32'b10111101001011100111010000110011 ;
        778: q <= 32'b10111101111100110001101011000101 ;
        779: q <= 32'b00111100010110010011001100110101 ;
        780: q <= 32'b00111101100111001110000100110110 ;
        781: q <= 32'b00111101001100100110011000101001 ;
        782: q <= 32'b00111101000010111011011010001100 ;
        783: q <= 32'b10111101100010100011101100101010 ;
        784: q <= 32'b10111100000111111110010100011010 ;
        785: q <= 32'b00111101001101011000001001100101 ;
        786: q <= 32'b10111110001010100001011100110100 ;
        787: q <= 32'b10111101100111010110101010011010 ;
        788: q <= 32'b10111011011010100011010101000111 ;
        789: q <= 32'b00111101000111000110110010111101 ;
        790: q <= 32'b00111101110101101110110101001111 ;
        791: q <= 32'b10111101111001110001110110000100 ;
        792: q <= 32'b00111110000000011001100111111000 ;
        793: q <= 32'b00111101100010011001000100110110 ;
        794: q <= 32'b10111101110101001001001101000100 ;
        795: q <= 32'b10111101100011110000101101101000 ;
        796: q <= 32'b00111101101100010010110011100010 ;
        797: q <= 32'b10111110000110101101011000000111 ;
        798: q <= 32'b10111010011001001001011010000111 ;
        799: q <= 32'b00111101000101100001100100111100 ;
        800: q <= 32'b10111100111101100011111001100110 ;
        801: q <= 32'b10111101001100111100111000000011 ;
        802: q <= 32'b10111100100111000001110010000000 ;
        803: q <= 32'b00111101110000101000111001110000 ;
        804: q <= 32'b10111101110001010100101001100101 ;
        805: q <= 32'b10111101110110101000000010010101 ;
        806: q <= 32'b00111101110011000000100011100000 ;
        807: q <= 32'b00111100100010001101001101110000 ;
        808: q <= 32'b00111100101100011111111011001110 ;
        809: q <= 32'b10111010110001001011010100001100 ;
        810: q <= 32'b10111100100000011100001110100001 ;
        811: q <= 32'b10111101101111110100000000101111 ;
        812: q <= 32'b10111101010001001110000001101000 ;
        813: q <= 32'b10111101100010110111111001110111 ;
        814: q <= 32'b10111101100010100001111100010010 ;
        815: q <= 32'b00111100101100101101000110101101 ;
        816: q <= 32'b10111100100000101001100001010000 ;
        817: q <= 32'b00111101110100110111101000010101 ;
        818: q <= 32'b00111101100011111011001100001100 ;
        819: q <= 32'b00111100011110010101101000110010 ;
        820: q <= 32'b00111100001000000001100111100011 ;
        821: q <= 32'b00111101101001010011100001110101 ;
        822: q <= 32'b10111101100011011010000000001111 ;
        823: q <= 32'b10111101100010010111101000000011 ;
        824: q <= 32'b10111011010010100001000111111100 ;
        825: q <= 32'b10111101010001101010101110101110 ;
        826: q <= 32'b00111100101111101110101000001111 ;
        827: q <= 32'b00111101001001001001101101101010 ;
        828: q <= 32'b00111101100001001100010000000111 ;
        829: q <= 32'b10111101001101100000101111001111 ;
        830: q <= 32'b00111011111011000100100101011101 ;
        831: q <= 32'b00111101101100110011001110110000 ;
        832: q <= 32'b10111100110011110101011101001110 ;
        833: q <= 32'b10111101010000010001100010100110 ;
        834: q <= 32'b00111101010111011001100100010100 ;
        835: q <= 32'b00111011101110111100100011110100 ;
        836: q <= 32'b00111011111001001110100111010011 ;
        837: q <= 32'b10111101100010010110111010101010 ;
        838: q <= 32'b10111101011001001101010100111110 ;
        839: q <= 32'b00111101010101010110001111001010 ;
        840: q <= 32'b10111100010101001010111101101010 ;
        841: q <= 32'b00111100001011000101100011000001 ;
        842: q <= 32'b10111101101101011010100101111011 ;
        843: q <= 32'b00111101101101011000101010101100 ;
        844: q <= 32'b00111100101000100001001000011010 ;
        845: q <= 32'b00111011010110011001011000101111 ;
        846: q <= 32'b10111101000100011110100011010000 ;
        847: q <= 32'b00111101111010010001001010100001 ;
        848: q <= 32'b00111101010110000010110101110001 ;
        849: q <= 32'b10111110000010101101111011011111 ;
        850: q <= 32'b10111110000011100010011100001000 ;
        851: q <= 32'b00111011100111001110110000001010 ;
        852: q <= 32'b10111101100011111110101101100000 ;
        853: q <= 32'b10111100111100000001101111100110 ;
        854: q <= 32'b00111011100110110101001000101010 ;
        855: q <= 32'b10111101100011100001010010110011 ;
        856: q <= 32'b10111101100001101110111000000111 ;
        857: q <= 32'b00111101100111011000110110000001 ;
        858: q <= 32'b10111101100011011011010010100100 ;
        859: q <= 32'b00111010011001110100111010011011 ;
        860: q <= 32'b00111110010000101101101010101000 ;
        861: q <= 32'b10111100110111000000111101011111 ;
        862: q <= 32'b00111011010001111110101011110100 ;
        863: q <= 32'b00111100111011000101100111111111 ;
        864: q <= 32'b10111101100110001011000110001011 ;
        865: q <= 32'b00111101001001011100101000000001 ;
        866: q <= 32'b00111101000101100011100110011100 ;
        867: q <= 32'b10111100011100100110010111011010 ;
        868: q <= 32'b10111101101011110110000100100110 ;
        869: q <= 32'b00111101110010111010001000100011 ;
        870: q <= 32'b10111101010110111101011110010011 ;
        871: q <= 32'b10111101100110110111000000111110 ;
        872: q <= 32'b00000000000000000000000000000000 ;
        873: q <= 32'b00000000000000000000000000000000 ;
        874: q <= 32'b00000000000000000000000000000000 ;
        875: q <= 32'b00000000000000000000000000000000 ;
        876: q <= 32'b00000000000000000000000000000000 ;
        877: q <= 32'b00000000000000000000000000000000 ;
        878: q <= 32'b00000000000000000000000000000000 ;
        879: q <= 32'b00000000000000000000000000000000 ;
        880: q <= 32'b00000000000000000000000000000000 ;
        881: q <= 32'b00000000000000000000000000000000 ;
        882: q <= 32'b00000000000000000000000000000000 ;
        883: q <= 32'b00000000000000000000000000000000 ;
        884: q <= 32'b00000000000000000000000000000000 ;
        885: q <= 32'b00000000000000000000000000000000 ;
        886: q <= 32'b00000000000000000000000000000000 ;
        887: q <= 32'b00000000000000000000000000000000 ;
        888: q <= 32'b00000000000000000000000000000000 ;
        889: q <= 32'b00000000000000000000000000000000 ;
        890: q <= 32'b00000000000000000000000000000000 ;
        891: q <= 32'b00000000000000000000000000000000 ;
        892: q <= 32'b00000000000000000000000000000000 ;
        893: q <= 32'b00000000000000000000000000000000 ;
        894: q <= 32'b00000000000000000000000000000000 ;
        895: q <= 32'b00000000000000000000000000000000 ;
        896: q <= 32'b10111101011101010101001011110001 ;
        897: q <= 32'b00111101100000111010000001001001 ;
        898: q <= 32'b00111101110010110110000101000011 ;
        899: q <= 32'b00111110000010110110010011100101 ;
        900: q <= 32'b00111101100110111101001101100100 ;
        901: q <= 32'b10111101111101100000011000011010 ;
        902: q <= 32'b00111101100111101110111000110110 ;
        903: q <= 32'b00111101111011111100110101011011 ;
        904: q <= 32'b10111110010000001010010110000001 ;
        905: q <= 32'b00111100001001111000111000001111 ;
        906: q <= 32'b10111101100001001000101110010111 ;
        907: q <= 32'b00111101100101111010100001000000 ;
        908: q <= 32'b00111101011011110111011010001100 ;
        909: q <= 32'b00111100000011101100100111100010 ;
        910: q <= 32'b10111101010111110001100010010010 ;
        911: q <= 32'b00111101100010110111001010100101 ;
        912: q <= 32'b00111101101000100000110101110000 ;
        913: q <= 32'b00111101000100110010001101101010 ;
        914: q <= 32'b00111101101100001000110001011110 ;
        915: q <= 32'b10111101011100011001100110100110 ;
        916: q <= 32'b00111100010011111000110010010000 ;
        917: q <= 32'b00111101111110110101101011001101 ;
        918: q <= 32'b10111101000011001101101011101001 ;
        919: q <= 32'b10111100001011001101010101001001 ;
        920: q <= 32'b10111101111010011000010000100001 ;
        921: q <= 32'b10111101010001000111000010101011 ;
        922: q <= 32'b00111101101010110010110000011000 ;
        923: q <= 32'b00111100101000011110100010111100 ;
        924: q <= 32'b10111101100100111101001011110010 ;
        925: q <= 32'b00111110001001110111001110010100 ;
        926: q <= 32'b00111101100001110110110100001001 ;
        927: q <= 32'b10111101001101001101111010110001 ;
        928: q <= 32'b10111101100110010011111100000101 ;
        929: q <= 32'b00111101100110101010111101110001 ;
        930: q <= 32'b10111110001000110000011100101011 ;
        931: q <= 32'b00111101101100011101011011000000 ;
        932: q <= 32'b10111100110101101101111010010110 ;
        933: q <= 32'b00111101010001111110111111101011 ;
        934: q <= 32'b00111101101011011110110010110010 ;
        935: q <= 32'b00111101001101100001111100111011 ;
        936: q <= 32'b00111101011010001111100000101110 ;
        937: q <= 32'b10111100110011100011111111110111 ;
        938: q <= 32'b10111101011010001101010100100010 ;
        939: q <= 32'b00111100100000001011011100000001 ;
        940: q <= 32'b00111100110111000010110110110110 ;
        941: q <= 32'b00111101100110000000011100010000 ;
        942: q <= 32'b10111100101100110001110101110111 ;
        943: q <= 32'b00111101010011010111101000111101 ;
        944: q <= 32'b10111101000001100011111010001101 ;
        945: q <= 32'b00111101011000100101001001110100 ;
        946: q <= 32'b00111101010000000000110011100101 ;
        947: q <= 32'b10111101110001111110110010110001 ;
        948: q <= 32'b00111100111010100011111001100010 ;
        949: q <= 32'b10111100101001001011011101011110 ;
        950: q <= 32'b10111100001111010001100101110000 ;
        951: q <= 32'b00111110000011001000101010011111 ;
        952: q <= 32'b00111011100001010100111000111100 ;
        953: q <= 32'b10111100101100000000110101001111 ;
        954: q <= 32'b10111101011101001011011101001111 ;
        955: q <= 32'b00111100101011100011100110010010 ;
        956: q <= 32'b10111101111110001110010100000000 ;
        957: q <= 32'b00111101001110100110111000101100 ;
        958: q <= 32'b10111010000001011001110011010001 ;
        959: q <= 32'b00111101011010011010011101110010 ;
        960: q <= 32'b10111100100101100111010100101101 ;
        961: q <= 32'b00111101010101100101101011100110 ;
        962: q <= 32'b00111110001011011000110011100000 ;
        963: q <= 32'b00111101100010110000011111010010 ;
        964: q <= 32'b00111101011011101001110001011011 ;
        965: q <= 32'b10111101010000101010101000100001 ;
        966: q <= 32'b10111101010000110010001111010011 ;
        967: q <= 32'b00111101100111010001111001000001 ;
        968: q <= 32'b00111011001100011111110100101010 ;
        969: q <= 32'b00111101111010101010011011000001 ;
        970: q <= 32'b10111100100110011010010110011100 ;
        971: q <= 32'b00111100011101110011001001010000 ;
        972: q <= 32'b00111101110111001100110111011100 ;
        973: q <= 32'b00111101011010001110100000100100 ;
        974: q <= 32'b10111110000001001100000110111010 ;
        975: q <= 32'b10111101011100001101110110110100 ;
        976: q <= 32'b00111110010100101000000000110100 ;
        977: q <= 32'b00111101000111011100010101001111 ;
        978: q <= 32'b00111110000000101101111010100000 ;
        979: q <= 32'b10111101011100101101001011001110 ;
        980: q <= 32'b10111100011100110111000001010110 ;
        981: q <= 32'b00111110000100101011111101001000 ;
        982: q <= 32'b10111101100011001001010111011101 ;
        983: q <= 32'b10111100000101111001110110010111 ;
        984: q <= 32'b10111100101011111111001101000101 ;
        985: q <= 32'b10111101110000011111101111011110 ;
        986: q <= 32'b00111100010010010011011100000101 ;
        987: q <= 32'b00111100110001101011011001101110 ;
        988: q <= 32'b00111101100011110100010011001010 ;
        989: q <= 32'b00111101111100010011101000010100 ;
        990: q <= 32'b00111100011011110111111100110010 ;
        991: q <= 32'b00111110010101101010011100010110 ;
        992: q <= 32'b10111101100011010010100010010000 ;
        993: q <= 32'b00111010001001101100000011100000 ;
        994: q <= 32'b00111110000100001111001001111100 ;
        995: q <= 32'b00111110000011101101000000100110 ;
        996: q <= 32'b10111101101010001110001100110011 ;
        997: q <= 32'b00111110000010111111001000100000 ;
        998: q <= 32'b10111101011001101100001100100011 ;
        999: q <= 32'b10111101100101010000011110001010 ;
        1000: q <= 32'b00000000000000000000000000000000 ;
        1001: q <= 32'b00000000000000000000000000000000 ;
        1002: q <= 32'b00000000000000000000000000000000 ;
        1003: q <= 32'b00000000000000000000000000000000 ;
        1004: q <= 32'b00000000000000000000000000000000 ;
        1005: q <= 32'b00000000000000000000000000000000 ;
        1006: q <= 32'b00000000000000000000000000000000 ;
        1007: q <= 32'b00000000000000000000000000000000 ;
        1008: q <= 32'b00000000000000000000000000000000 ;
        1009: q <= 32'b00000000000000000000000000000000 ;
        1010: q <= 32'b00000000000000000000000000000000 ;
        1011: q <= 32'b00000000000000000000000000000000 ;
        1012: q <= 32'b00000000000000000000000000000000 ;
        1013: q <= 32'b00000000000000000000000000000000 ;
        1014: q <= 32'b00000000000000000000000000000000 ;
        1015: q <= 32'b00000000000000000000000000000000 ;
        1016: q <= 32'b00000000000000000000000000000000 ;
        1017: q <= 32'b00000000000000000000000000000000 ;
        1018: q <= 32'b00000000000000000000000000000000 ;
        1019: q <= 32'b00000000000000000000000000000000 ;
        1020: q <= 32'b00000000000000000000000000000000 ;
        1021: q <= 32'b00000000000000000000000000000000 ;
        1022: q <= 32'b00000000000000000000000000000000 ;
        1023: q <= 32'b00000000000000000000000000000000 ;
        1024: q <= 32'b00111100100011111110001110100110 ;
        1025: q <= 32'b10111101010000010010100101110001 ;
        1026: q <= 32'b10111101000010000110001011110001 ;
        1027: q <= 32'b10111101110100100111001010111101 ;
        1028: q <= 32'b10111101000100001010110000010100 ;
        1029: q <= 32'b00111101100111011010110110000101 ;
        1030: q <= 32'b10111101001110100001001010110010 ;
        1031: q <= 32'b00111101011101010101111010100100 ;
        1032: q <= 32'b10111100111110110111010010000011 ;
        1033: q <= 32'b00111011100000100010001001001011 ;
        1034: q <= 32'b00111101101001100111100101111011 ;
        1035: q <= 32'b10111101011001100000000111010101 ;
        1036: q <= 32'b10111101011010010110010010101000 ;
        1037: q <= 32'b10111101100100110110010100101001 ;
        1038: q <= 32'b00111101100011110000011110101001 ;
        1039: q <= 32'b10111110000000010001110011111110 ;
        1040: q <= 32'b10111101100101101101110100010110 ;
        1041: q <= 32'b10111101100101001000111110010101 ;
        1042: q <= 32'b00111101101110010011011001110000 ;
        1043: q <= 32'b10111101101000101100010000111111 ;
        1044: q <= 32'b00111011110001111011000101111111 ;
        1045: q <= 32'b10111100111100101000011011101001 ;
        1046: q <= 32'b00111011100011101101100100010101 ;
        1047: q <= 32'b00111101100111001111001101110100 ;
        1048: q <= 32'b10111101101111000100111011011111 ;
        1049: q <= 32'b00111101100111110111000000111000 ;
        1050: q <= 32'b10111101111110000001110011010001 ;
        1051: q <= 32'b10111011001111010010110101111111 ;
        1052: q <= 32'b10111101000110110110011001011000 ;
        1053: q <= 32'b00111101001010001000111001101110 ;
        1054: q <= 32'b00111101000101101011100000001100 ;
        1055: q <= 32'b10111101110011100010111000111000 ;
        1056: q <= 32'b10111101101100001101100101010001 ;
        1057: q <= 32'b00111100100101001110011000011110 ;
        1058: q <= 32'b00111101001100110010000011111011 ;
        1059: q <= 32'b10111101100010011000111111110101 ;
        1060: q <= 32'b10111101100000111100011100000101 ;
        1061: q <= 32'b00111100000011010110100101010010 ;
        1062: q <= 32'b00111100001011110111111101100000 ;
        1063: q <= 32'b10111010101010110000001000110001 ;
        1064: q <= 32'b10111011101000011100010001011110 ;
        1065: q <= 32'b10111101011100000110010000111000 ;
        1066: q <= 32'b00111101011001101011110111111001 ;
        1067: q <= 32'b10111101101110101101000111100000 ;
        1068: q <= 32'b00111101100001011000011110100010 ;
        1069: q <= 32'b10111101110010000101010011001110 ;
        1070: q <= 32'b10111100001001010101001001101111 ;
        1071: q <= 32'b00111101100011110111010101000111 ;
        1072: q <= 32'b10111101110101001100000011001001 ;
        1073: q <= 32'b00111100111110111011000010000000 ;
        1074: q <= 32'b00111101101011010101110010111111 ;
        1075: q <= 32'b10111101101101010001001101000001 ;
        1076: q <= 32'b10111101100011101111001101011001 ;
        1077: q <= 32'b10111101100001000110110111110101 ;
        1078: q <= 32'b10111101110000000111100101011101 ;
        1079: q <= 32'b10111011001100001000110010001000 ;
        1080: q <= 32'b00111100110010110110101111001011 ;
        1081: q <= 32'b10111101010110111111100100100101 ;
        1082: q <= 32'b10111101010001001000000110000000 ;
        1083: q <= 32'b10111101001001000010110111101110 ;
        1084: q <= 32'b00111100111110110111010100010011 ;
        1085: q <= 32'b00111101011111101000100100010110 ;
        1086: q <= 32'b00111101101011101100100000111110 ;
        1087: q <= 32'b00111011001001001010111111001001 ;
        1088: q <= 32'b00111101000100011001101010011000 ;
        1089: q <= 32'b10111101010011001000110011011110 ;
        1090: q <= 32'b00111101010100111100110111010011 ;
        1091: q <= 32'b10111101100010011000110100010111 ;
        1092: q <= 32'b10111101000111000110010000110111 ;
        1093: q <= 32'b10111100001011111101101111100101 ;
        1094: q <= 32'b10111101100011110001001010011100 ;
        1095: q <= 32'b10111101101010001011010101001101 ;
        1096: q <= 32'b00111100000110101101111110111010 ;
        1097: q <= 32'b00111100111110000011101111101100 ;
        1098: q <= 32'b10111101010001011110110000101101 ;
        1099: q <= 32'b10111101001001100100100101111001 ;
        1100: q <= 32'b10111100101011100010100000010001 ;
        1101: q <= 32'b10111101110011111110111011100000 ;
        1102: q <= 32'b10111101011111011000011100000111 ;
        1103: q <= 32'b10111100110010011110110110111000 ;
        1104: q <= 32'b00111100110010010110011000111101 ;
        1105: q <= 32'b10111101100001110100011101010010 ;
        1106: q <= 32'b10111101010111010110100001111010 ;
        1107: q <= 32'b10111101011101100011100110000101 ;
        1108: q <= 32'b00111101011000010100101011111001 ;
        1109: q <= 32'b00111101100000010011011110101101 ;
        1110: q <= 32'b00111101100010111111100010100001 ;
        1111: q <= 32'b00111101101000111001101111010100 ;
        1112: q <= 32'b00111011100011111100110001111100 ;
        1113: q <= 32'b00111101001100111000111111010011 ;
        1114: q <= 32'b00111011000110011101000010100001 ;
        1115: q <= 32'b00111101011011001101101011011011 ;
        1116: q <= 32'b00111101011110100001010101101111 ;
        1117: q <= 32'b10111100111000000110111000010000 ;
        1118: q <= 32'b00111010001110011111101111011100 ;
        1119: q <= 32'b10111100101001110110000000110110 ;
        1120: q <= 32'b10111101110010010010001110110111 ;
        1121: q <= 32'b10111100110010011110101010111010 ;
        1122: q <= 32'b10111101100001101100111110110010 ;
        1123: q <= 32'b00111101001000100101100110100111 ;
        1124: q <= 32'b00111101010100100010011000010101 ;
        1125: q <= 32'b10111010000000100011100100010001 ;
        1126: q <= 32'b10111101100001111111001010000000 ;
        1127: q <= 32'b10111101010100001001100101110111 ;
        1128: q <= 32'b00000000000000000000000000000000 ;
        1129: q <= 32'b00000000000000000000000000000000 ;
        1130: q <= 32'b00000000000000000000000000000000 ;
        1131: q <= 32'b00000000000000000000000000000000 ;
        1132: q <= 32'b00000000000000000000000000000000 ;
        1133: q <= 32'b00000000000000000000000000000000 ;
        1134: q <= 32'b00000000000000000000000000000000 ;
        1135: q <= 32'b00000000000000000000000000000000 ;
        1136: q <= 32'b00000000000000000000000000000000 ;
        1137: q <= 32'b00000000000000000000000000000000 ;
        1138: q <= 32'b00000000000000000000000000000000 ;
        1139: q <= 32'b00000000000000000000000000000000 ;
        1140: q <= 32'b00000000000000000000000000000000 ;
        1141: q <= 32'b00000000000000000000000000000000 ;
        1142: q <= 32'b00000000000000000000000000000000 ;
        1143: q <= 32'b00000000000000000000000000000000 ;
        1144: q <= 32'b00000000000000000000000000000000 ;
        1145: q <= 32'b00000000000000000000000000000000 ;
        1146: q <= 32'b00000000000000000000000000000000 ;
        1147: q <= 32'b00000000000000000000000000000000 ;
        1148: q <= 32'b00000000000000000000000000000000 ;
        1149: q <= 32'b00000000000000000000000000000000 ;
        1150: q <= 32'b00000000000000000000000000000000 ;
        1151: q <= 32'b00000000000000000000000000000000 ;
        1152: q <= 32'b10111100110101100100111010010111 ;
        1153: q <= 32'b00111110001110010001101001010011 ;
        1154: q <= 32'b10111100100111111000101110000000 ;
        1155: q <= 32'b10111100110111101000111110001001 ;
        1156: q <= 32'b00111101101000100110110001101011 ;
        1157: q <= 32'b00111101001000111000111000001101 ;
        1158: q <= 32'b10111101000010001101100101001100 ;
        1159: q <= 32'b10111101001001010011010001000000 ;
        1160: q <= 32'b00111101100001100111101011100001 ;
        1161: q <= 32'b00111101001010000001001011110000 ;
        1162: q <= 32'b10111101100000100010111010011011 ;
        1163: q <= 32'b10111101100011110100010100010010 ;
        1164: q <= 32'b00111100100111000011011110011100 ;
        1165: q <= 32'b10111101110100011101011110000001 ;
        1166: q <= 32'b10111101101000001011100100000101 ;
        1167: q <= 32'b00111100000010100001111101001000 ;
        1168: q <= 32'b00111101111101000000011111000111 ;
        1169: q <= 32'b00111100101010010010001101101001 ;
        1170: q <= 32'b00111110001011000111011111101101 ;
        1171: q <= 32'b00111101000000000101001110101110 ;
        1172: q <= 32'b10111101110101111111011101000100 ;
        1173: q <= 32'b10111101000000011001000001101001 ;
        1174: q <= 32'b10111101110001101011100110010000 ;
        1175: q <= 32'b10111101101011100111110000111110 ;
        1176: q <= 32'b10111100110010101011010001000110 ;
        1177: q <= 32'b10111101101001110011010000101001 ;
        1178: q <= 32'b10111110000001111011011001101101 ;
        1179: q <= 32'b00111100100110000011100010110100 ;
        1180: q <= 32'b00111101010110011010010110111000 ;
        1181: q <= 32'b00111101110110111001011010111101 ;
        1182: q <= 32'b00111101111000100011001011010001 ;
        1183: q <= 32'b00111101100010001011101000110111 ;
        1184: q <= 32'b00111100110111100100110010011100 ;
        1185: q <= 32'b00111100110111101000000111101010 ;
        1186: q <= 32'b10111101010001011001101101011010 ;
        1187: q <= 32'b00111101110000100111000010111010 ;
        1188: q <= 32'b00111101000110010101011111000111 ;
        1189: q <= 32'b10111101001000011100010001111100 ;
        1190: q <= 32'b10111101110000011101100100011000 ;
        1191: q <= 32'b00111101000010100011101101010011 ;
        1192: q <= 32'b00111101100000110110000110100000 ;
        1193: q <= 32'b10111011111100010111001001001111 ;
        1194: q <= 32'b00111100111010011011000011111010 ;
        1195: q <= 32'b00111101100010100100110110000011 ;
        1196: q <= 32'b10111101110010101111110111000011 ;
        1197: q <= 32'b10111101101101010100001100000101 ;
        1198: q <= 32'b00111100001010100100110101000010 ;
        1199: q <= 32'b10111101100011010001001101000110 ;
        1200: q <= 32'b00111100010110011000000011111000 ;
        1201: q <= 32'b10111100011100000011000000011000 ;
        1202: q <= 32'b10111101010001010101000110000000 ;
        1203: q <= 32'b00111101101101010001001001001111 ;
        1204: q <= 32'b10111101110000010101000000111000 ;
        1205: q <= 32'b00111101010011100100011111000010 ;
        1206: q <= 32'b10111101010101100010011010111001 ;
        1207: q <= 32'b10111101001001001011111011110011 ;
        1208: q <= 32'b10111101010100100101010111110010 ;
        1209: q <= 32'b10111101101111110111110111000100 ;
        1210: q <= 32'b10111100000001111000111011101101 ;
        1211: q <= 32'b10111100000110111100111011101101 ;
        1212: q <= 32'b00111101010000100110011011101101 ;
        1213: q <= 32'b10111101110000110100011000100011 ;
        1214: q <= 32'b10111100101110001100001000100010 ;
        1215: q <= 32'b00111101010110001011101111100000 ;
        1216: q <= 32'b10111101011111011000111111111010 ;
        1217: q <= 32'b10111101110010001010001001010100 ;
        1218: q <= 32'b10111100111010110111101110110011 ;
        1219: q <= 32'b00111100101101101000011100101010 ;
        1220: q <= 32'b10111011111011000100000111111011 ;
        1221: q <= 32'b00111101101111011000110010101110 ;
        1222: q <= 32'b00111101110000011111011001110101 ;
        1223: q <= 32'b00111101110001000011001100110111 ;
        1224: q <= 32'b00111101110011001101001000001011 ;
        1225: q <= 32'b10111101100011001110010110100110 ;
        1226: q <= 32'b00111101010110111010010001111110 ;
        1227: q <= 32'b00111110000011101110100010111010 ;
        1228: q <= 32'b10111101101110110011100000001100 ;
        1229: q <= 32'b00111101001011101100110000100111 ;
        1230: q <= 32'b10111101000010100111100110110110 ;
        1231: q <= 32'b00111100000101101000010000111111 ;
        1232: q <= 32'b00111101100100001000011100101001 ;
        1233: q <= 32'b10111100001000011100101000101101 ;
        1234: q <= 32'b00111101001100000101100010100001 ;
        1235: q <= 32'b00111101100001101010010111001000 ;
        1236: q <= 32'b00111100011101111000110011101111 ;
        1237: q <= 32'b00111101001000101010011000010000 ;
        1238: q <= 32'b00111101100010101100011100101110 ;
        1239: q <= 32'b10111101000000111111111001000110 ;
        1240: q <= 32'b00111101001111110101011101001001 ;
        1241: q <= 32'b10111101010010010010111101101100 ;
        1242: q <= 32'b00111101101000100011110011010000 ;
        1243: q <= 32'b00111101100001001110011100110100 ;
        1244: q <= 32'b10111110001010100001100011010011 ;
        1245: q <= 32'b10111100100011100010001111101000 ;
        1246: q <= 32'b00111101110011010101001001100101 ;
        1247: q <= 32'b10111101001010000100110010100110 ;
        1248: q <= 32'b00111101110110011010111100111001 ;
        1249: q <= 32'b00111011101101001000110000000111 ;
        1250: q <= 32'b00111101101110100100001110001100 ;
        1251: q <= 32'b00111110001100110110011100010111 ;
        1252: q <= 32'b00111101101110011000010000001011 ;
        1253: q <= 32'b10111101010001110010011101011010 ;
        1254: q <= 32'b00111100100011110011011000100101 ;
        1255: q <= 32'b00111101000010110010101101100111 ;
        1256: q <= 32'b00000000000000000000000000000000 ;
        1257: q <= 32'b00000000000000000000000000000000 ;
        1258: q <= 32'b00000000000000000000000000000000 ;
        1259: q <= 32'b00000000000000000000000000000000 ;
        1260: q <= 32'b00000000000000000000000000000000 ;
        1261: q <= 32'b00000000000000000000000000000000 ;
        1262: q <= 32'b00000000000000000000000000000000 ;
        1263: q <= 32'b00000000000000000000000000000000 ;
        1264: q <= 32'b00000000000000000000000000000000 ;
        1265: q <= 32'b00000000000000000000000000000000 ;
        1266: q <= 32'b00000000000000000000000000000000 ;
        1267: q <= 32'b00000000000000000000000000000000 ;
        1268: q <= 32'b00000000000000000000000000000000 ;
        1269: q <= 32'b00000000000000000000000000000000 ;
        1270: q <= 32'b00000000000000000000000000000000 ;
        1271: q <= 32'b00000000000000000000000000000000 ;
        1272: q <= 32'b00000000000000000000000000000000 ;
        1273: q <= 32'b00000000000000000000000000000000 ;
        1274: q <= 32'b00000000000000000000000000000000 ;
        1275: q <= 32'b00000000000000000000000000000000 ;
        1276: q <= 32'b00000000000000000000000000000000 ;
        1277: q <= 32'b00000000000000000000000000000000 ;
        1278: q <= 32'b00000000000000000000000000000000 ;
        1279: q <= 32'b00000000000000000000000000000000 ;
        1280: q <= 32'b00111110000110001111001001111001 ;
        1281: q <= 32'b00111101111011001101110011011010 ;
        1282: q <= 32'b00111101110010011011111010100100 ;
        1283: q <= 32'b10111100110101001000011011001001 ;
        1284: q <= 32'b00111101001101010111000011110001 ;
        1285: q <= 32'b00111010100000110010000001000011 ;
        1286: q <= 32'b00111101011000101010101111100011 ;
        1287: q <= 32'b00111101100010011111100001011111 ;
        1288: q <= 32'b10111101100010000000011010100111 ;
        1289: q <= 32'b00111010101101000111011100011111 ;
        1290: q <= 32'b10111100001011111010111000100010 ;
        1291: q <= 32'b00111101001110111101111101111010 ;
        1292: q <= 32'b10111101001110111111100010110001 ;
        1293: q <= 32'b10111101011110001101100010111101 ;
        1294: q <= 32'b10111101100010100001110010110010 ;
        1295: q <= 32'b10111101100010000111101000111110 ;
        1296: q <= 32'b00111011111001010100010000010100 ;
        1297: q <= 32'b10111100110101110101001110001101 ;
        1298: q <= 32'b10111101010100001111010101111100 ;
        1299: q <= 32'b10111101010000111101111101010000 ;
        1300: q <= 32'b10111101100101101000000100001000 ;
        1301: q <= 32'b10111101000000001100011100101100 ;
        1302: q <= 32'b00111101001000110011111001001100 ;
        1303: q <= 32'b00111101000100101000110110000101 ;
        1304: q <= 32'b10111100001110001010000010011000 ;
        1305: q <= 32'b10111100100110011011001010011100 ;
        1306: q <= 32'b00111100001111100101111001010011 ;
        1307: q <= 32'b10111011101011100001111011001110 ;
        1308: q <= 32'b10111101011001001110011110111100 ;
        1309: q <= 32'b00111101100011111110101101110101 ;
        1310: q <= 32'b10111101010100001110011000011010 ;
        1311: q <= 32'b10111101011011000111100111011000 ;
        1312: q <= 32'b00111101110101100110110000101010 ;
        1313: q <= 32'b00111101010001010000000000111100 ;
        1314: q <= 32'b10111101101011011000000110100001 ;
        1315: q <= 32'b00111101101110000111101111110111 ;
        1316: q <= 32'b10111101100110110010101001011111 ;
        1317: q <= 32'b10111011011010100110010110010010 ;
        1318: q <= 32'b00111100101111111010100001100111 ;
        1319: q <= 32'b00111100110011000111010001010110 ;
        1320: q <= 32'b00111101010110010010101111001001 ;
        1321: q <= 32'b10111010110000111011000010101101 ;
        1322: q <= 32'b10111101001000011000010010010100 ;
        1323: q <= 32'b00111101100110001010110101010001 ;
        1324: q <= 32'b10111100100100101001110100001110 ;
        1325: q <= 32'b10111001110111011010011001011110 ;
        1326: q <= 32'b00111101110001010100101000111100 ;
        1327: q <= 32'b10111101011011110100001000011010 ;
        1328: q <= 32'b00111100110111000111010011100111 ;
        1329: q <= 32'b10111101001101101101000000010110 ;
        1330: q <= 32'b10111101100011011110110001110101 ;
        1331: q <= 32'b10111101010110110110000011111000 ;
        1332: q <= 32'b00111100110000011000010000011010 ;
        1333: q <= 32'b00111101101001001001101110111010 ;
        1334: q <= 32'b00111101011110111110110000000100 ;
        1335: q <= 32'b10111101100100110010000110010101 ;
        1336: q <= 32'b10111101100110101111010111010111 ;
        1337: q <= 32'b10111101000011111010110110001100 ;
        1338: q <= 32'b10111101100010000011000111000100 ;
        1339: q <= 32'b00111101010000000000010010101100 ;
        1340: q <= 32'b10111101100001001110001001011011 ;
        1341: q <= 32'b00111100101011011101100110001011 ;
        1342: q <= 32'b00111101011000001110110101011101 ;
        1343: q <= 32'b00111101100010100000001101110001 ;
        1344: q <= 32'b10111100110011100011110001111111 ;
        1345: q <= 32'b10111000010101100111010010010110 ;
        1346: q <= 32'b00111100101111001100110000110010 ;
        1347: q <= 32'b10111101001001100001000101001111 ;
        1348: q <= 32'b10111101010100100001000100111110 ;
        1349: q <= 32'b00111100100010011011010001001110 ;
        1350: q <= 32'b00111101101001000101011011011011 ;
        1351: q <= 32'b10111100101111011011010110000100 ;
        1352: q <= 32'b10111100111100101101000110111110 ;
        1353: q <= 32'b10111101001011110101011100101011 ;
        1354: q <= 32'b00111101110101001110101110010011 ;
        1355: q <= 32'b00111100011101000100011011110011 ;
        1356: q <= 32'b10111101101100010001101000011100 ;
        1357: q <= 32'b00111101011010111100001001100110 ;
        1358: q <= 32'b00111101101111010101101111000110 ;
        1359: q <= 32'b10111101101000111001010101011010 ;
        1360: q <= 32'b00111101101110100110000010000001 ;
        1361: q <= 32'b10111100110111001011110111101100 ;
        1362: q <= 32'b00111101101011110010011010100111 ;
        1363: q <= 32'b00111101001110111000111000001011 ;
        1364: q <= 32'b10111101101100100100100101011100 ;
        1365: q <= 32'b10111101010010011010000001010000 ;
        1366: q <= 32'b00111101100111010111000100010001 ;
        1367: q <= 32'b00111101100110000011111101001111 ;
        1368: q <= 32'b00111100101010001111110111110101 ;
        1369: q <= 32'b00111101101010001001111000101011 ;
        1370: q <= 32'b00111101101000100010000001000101 ;
        1371: q <= 32'b10111100100001000001111001010001 ;
        1372: q <= 32'b10111101100001111000100000100111 ;
        1373: q <= 32'b10111101001100110000010001010000 ;
        1374: q <= 32'b10111101100110000110110011001011 ;
        1375: q <= 32'b00111101010110101101110100111110 ;
        1376: q <= 32'b00111101101010000101001000100010 ;
        1377: q <= 32'b10111101010101001110000000000101 ;
        1378: q <= 32'b00111101001111010000101010011100 ;
        1379: q <= 32'b10111100110111011110010000010001 ;
        1380: q <= 32'b00111101000000101101010000111111 ;
        1381: q <= 32'b10111101000100100101101111010100 ;
        1382: q <= 32'b00111101101001101010001010011111 ;
        1383: q <= 32'b00111101110101100011011111010101 ;
        1384: q <= 32'b00000000000000000000000000000000 ;
        1385: q <= 32'b00000000000000000000000000000000 ;
        1386: q <= 32'b00000000000000000000000000000000 ;
        1387: q <= 32'b00000000000000000000000000000000 ;
        1388: q <= 32'b00000000000000000000000000000000 ;
        1389: q <= 32'b00000000000000000000000000000000 ;
        1390: q <= 32'b00000000000000000000000000000000 ;
        1391: q <= 32'b00000000000000000000000000000000 ;
        1392: q <= 32'b00000000000000000000000000000000 ;
        1393: q <= 32'b00000000000000000000000000000000 ;
        1394: q <= 32'b00000000000000000000000000000000 ;
        1395: q <= 32'b00000000000000000000000000000000 ;
        1396: q <= 32'b00000000000000000000000000000000 ;
        1397: q <= 32'b00000000000000000000000000000000 ;
        1398: q <= 32'b00000000000000000000000000000000 ;
        1399: q <= 32'b00000000000000000000000000000000 ;
        1400: q <= 32'b00000000000000000000000000000000 ;
        1401: q <= 32'b00000000000000000000000000000000 ;
        1402: q <= 32'b00000000000000000000000000000000 ;
        1403: q <= 32'b00000000000000000000000000000000 ;
        1404: q <= 32'b00000000000000000000000000000000 ;
        1405: q <= 32'b00000000000000000000000000000000 ;
        1406: q <= 32'b00000000000000000000000000000000 ;
        1407: q <= 32'b00000000000000000000000000000000 ;
        1408: q <= 32'b00111011101100010111001100101101 ;
        1409: q <= 32'b10111110000110110100010110011111 ;
        1410: q <= 32'b10111100000110100001111111011001 ;
        1411: q <= 32'b00111101110010011011001010001111 ;
        1412: q <= 32'b10111101000001100111010101111000 ;
        1413: q <= 32'b10111101001011111111001110011011 ;
        1414: q <= 32'b10111101100100110001100100110100 ;
        1415: q <= 32'b00111101000101111110110101100111 ;
        1416: q <= 32'b10111101111100100101101000001011 ;
        1417: q <= 32'b00111101101101010011111110000110 ;
        1418: q <= 32'b10111101111010100001110000001101 ;
        1419: q <= 32'b10111101111101010001100110111101 ;
        1420: q <= 32'b00111101100000110010101100111110 ;
        1421: q <= 32'b00111011111101111111010110111100 ;
        1422: q <= 32'b10111011100110001010000001010011 ;
        1423: q <= 32'b10111101101111010110011101000000 ;
        1424: q <= 32'b10111101110010010000001011100000 ;
        1425: q <= 32'b00111101110000110011001101101011 ;
        1426: q <= 32'b10111101100111111010111101000101 ;
        1427: q <= 32'b00111110000000111100110001011011 ;
        1428: q <= 32'b10111101010010010111111000010010 ;
        1429: q <= 32'b00111101111111001000001110101011 ;
        1430: q <= 32'b10111101101010011001111000100001 ;
        1431: q <= 32'b10111011010111110001101000010011 ;
        1432: q <= 32'b10111100011110111001011110001001 ;
        1433: q <= 32'b00111101010010101001111101101100 ;
        1434: q <= 32'b10111101010000111011000111101110 ;
        1435: q <= 32'b10111101010111111101110001101110 ;
        1436: q <= 32'b00111110001011010010000111110010 ;
        1437: q <= 32'b00111100111100101111000111101010 ;
        1438: q <= 32'b00111110000110011100011101100000 ;
        1439: q <= 32'b00111101001010001000010100100101 ;
        1440: q <= 32'b00111011001001010001001111100111 ;
        1441: q <= 32'b00111101000000010010010101001001 ;
        1442: q <= 32'b10111101111100010011110001110100 ;
        1443: q <= 32'b00111101101111110001100010111001 ;
        1444: q <= 32'b00111101100100000111110110101001 ;
        1445: q <= 32'b10111101000111001110010000001000 ;
        1446: q <= 32'b00111101110101101011000001000101 ;
        1447: q <= 32'b00111101110110101011010001101000 ;
        1448: q <= 32'b10111110001010100000010000000000 ;
        1449: q <= 32'b10111101101010111000001110111000 ;
        1450: q <= 32'b00111010101010010010001111010100 ;
        1451: q <= 32'b00111101111110111100000000100001 ;
        1452: q <= 32'b10111101101100001100111010110010 ;
        1453: q <= 32'b00111101110000101110000001100000 ;
        1454: q <= 32'b10111101100000000011100100101110 ;
        1455: q <= 32'b00111100000110101001101000111011 ;
        1456: q <= 32'b10111101100010111100000100011111 ;
        1457: q <= 32'b00111101001100001101001001111110 ;
        1458: q <= 32'b00111101110011100111100110000011 ;
        1459: q <= 32'b00111100110111101001101110101110 ;
        1460: q <= 32'b00111010100111000001111110010011 ;
        1461: q <= 32'b10111100010100010100101010011100 ;
        1462: q <= 32'b00111101111010010101001100111001 ;
        1463: q <= 32'b10111010101000101111010010101011 ;
        1464: q <= 32'b00111101100000111111110011000110 ;
        1465: q <= 32'b00111101011011011011100111110111 ;
        1466: q <= 32'b10111110000000111001000010010010 ;
        1467: q <= 32'b10111101000000100100100001000101 ;
        1468: q <= 32'b10111101011111110100110000111010 ;
        1469: q <= 32'b00111101110100001000010110000000 ;
        1470: q <= 32'b10111100101010011010111101100001 ;
        1471: q <= 32'b00111101101000001101011101111011 ;
        1472: q <= 32'b00111101001110010101001010100000 ;
        1473: q <= 32'b00111101000111100000110101011110 ;
        1474: q <= 32'b10111101010001001000110110001110 ;
        1475: q <= 32'b10111101010010111110110001001101 ;
        1476: q <= 32'b00111100100110010001101110011001 ;
        1477: q <= 32'b00111101110100100100111011110011 ;
        1478: q <= 32'b10111100000000000010101001111011 ;
        1479: q <= 32'b10111110001100011000101101011111 ;
        1480: q <= 32'b10111101101100001101010001001100 ;
        1481: q <= 32'b00111101111101000101110110010001 ;
        1482: q <= 32'b10111100110101001011100110101111 ;
        1483: q <= 32'b00111100110001110011010010111110 ;
        1484: q <= 32'b10111100111110001010101100010111 ;
        1485: q <= 32'b10111101100110111010101110100011 ;
        1486: q <= 32'b00111110000100010011111000000010 ;
        1487: q <= 32'b00111100101000111100101010001100 ;
        1488: q <= 32'b10111011111101100100011010110001 ;
        1489: q <= 32'b00111100100000010000000111011011 ;
        1490: q <= 32'b00111110100100010111110111101100 ;
        1491: q <= 32'b00111101111100100100111111110100 ;
        1492: q <= 32'b00111100001100110001001101100100 ;
        1493: q <= 32'b10111100110011110001001010110100 ;
        1494: q <= 32'b00111011010011010101100011010010 ;
        1495: q <= 32'b00111101101100010010110101100111 ;
        1496: q <= 32'b10111011110101001001110011011110 ;
        1497: q <= 32'b10111100111110100110001011001110 ;
        1498: q <= 32'b10111101010111010000000100110011 ;
        1499: q <= 32'b00111101010111100111110011101110 ;
        1500: q <= 32'b00111100110110000111010011100001 ;
        1501: q <= 32'b00111100101000011001001001001000 ;
        1502: q <= 32'b10111100111001001000110001010010 ;
        1503: q <= 32'b00111101000100001010011101110101 ;
        1504: q <= 32'b00111110000001001011110101001001 ;
        1505: q <= 32'b10111101011101110001110000101010 ;
        1506: q <= 32'b10111101111000111000111100010000 ;
        1507: q <= 32'b00111110000001101000001100111000 ;
        1508: q <= 32'b00111101110100000110111111010010 ;
        1509: q <= 32'b00111110000000101111110001000110 ;
        1510: q <= 32'b00111101101100110110000011100000 ;
        1511: q <= 32'b00111101100011011011001110010110 ;
        1512: q <= 32'b00000000000000000000000000000000 ;
        1513: q <= 32'b00000000000000000000000000000000 ;
        1514: q <= 32'b00000000000000000000000000000000 ;
        1515: q <= 32'b00000000000000000000000000000000 ;
        1516: q <= 32'b00000000000000000000000000000000 ;
        1517: q <= 32'b00000000000000000000000000000000 ;
        1518: q <= 32'b00000000000000000000000000000000 ;
        1519: q <= 32'b00000000000000000000000000000000 ;
        1520: q <= 32'b00000000000000000000000000000000 ;
        1521: q <= 32'b00000000000000000000000000000000 ;
        1522: q <= 32'b00000000000000000000000000000000 ;
        1523: q <= 32'b00000000000000000000000000000000 ;
        1524: q <= 32'b00000000000000000000000000000000 ;
        1525: q <= 32'b00000000000000000000000000000000 ;
        1526: q <= 32'b00000000000000000000000000000000 ;
        1527: q <= 32'b00000000000000000000000000000000 ;
        1528: q <= 32'b00000000000000000000000000000000 ;
        1529: q <= 32'b00000000000000000000000000000000 ;
        1530: q <= 32'b00000000000000000000000000000000 ;
        1531: q <= 32'b00000000000000000000000000000000 ;
        1532: q <= 32'b00000000000000000000000000000000 ;
        1533: q <= 32'b00000000000000000000000000000000 ;
        1534: q <= 32'b00000000000000000000000000000000 ;
        1535: q <= 32'b00000000000000000000000000000000 ;
        1536: q <= 32'b10111101100010101010101000100001 ;
        1537: q <= 32'b00111101101101010001100010001011 ;
        1538: q <= 32'b00111101101010001000110001110001 ;
        1539: q <= 32'b10111101101101101110101111011010 ;
        1540: q <= 32'b10111101100111100100110111001110 ;
        1541: q <= 32'b10111100011110000100110101010100 ;
        1542: q <= 32'b10111101110111011100101101110101 ;
        1543: q <= 32'b10111101101100111000100110011011 ;
        1544: q <= 32'b10111100011111101011000101111011 ;
        1545: q <= 32'b10111101101001101100111000000001 ;
        1546: q <= 32'b10111101001110001101011001100101 ;
        1547: q <= 32'b10111101000001001110101100011010 ;
        1548: q <= 32'b00111100000111001111110100010000 ;
        1549: q <= 32'b00111101011011001011111111011000 ;
        1550: q <= 32'b10111101010000011010010101101000 ;
        1551: q <= 32'b10111101011101000110001011111010 ;
        1552: q <= 32'b00111101100111110010111111001010 ;
        1553: q <= 32'b00111110010001110000001000000001 ;
        1554: q <= 32'b10111100001001010001010011111100 ;
        1555: q <= 32'b10111110001010100111101100100100 ;
        1556: q <= 32'b10111100000101110100100111110101 ;
        1557: q <= 32'b10111110000111010111110111011001 ;
        1558: q <= 32'b00111110001010111110011000111100 ;
        1559: q <= 32'b00111101111010010100000111101111 ;
        1560: q <= 32'b10111100111100100110101000110010 ;
        1561: q <= 32'b10111101110000101101110100010110 ;
        1562: q <= 32'b10111101111100010011010111110001 ;
        1563: q <= 32'b00111101100001110101111010001011 ;
        1564: q <= 32'b00111101000001111000011111010110 ;
        1565: q <= 32'b00111101011011010100111101100100 ;
        1566: q <= 32'b00111100100110001101101000011010 ;
        1567: q <= 32'b00111101010110111010000111101111 ;
        1568: q <= 32'b10111101111100111001100111100111 ;
        1569: q <= 32'b10111101110010100001000010111111 ;
        1570: q <= 32'b10111110000101010110010111111010 ;
        1571: q <= 32'b10111101001001111111110100110011 ;
        1572: q <= 32'b00111101110101111100101011111011 ;
        1573: q <= 32'b10111101100111010111100111011111 ;
        1574: q <= 32'b00111100011101110111100011010111 ;
        1575: q <= 32'b10111100101101001010110011111010 ;
        1576: q <= 32'b10111101011001111111100000100011 ;
        1577: q <= 32'b00111100111001100000011110001100 ;
        1578: q <= 32'b10111101000100001010110100001100 ;
        1579: q <= 32'b00111101101010110101111001000011 ;
        1580: q <= 32'b10111101000110011111010011001011 ;
        1581: q <= 32'b10111011001000011111011110011001 ;
        1582: q <= 32'b10111101101001111110100000101111 ;
        1583: q <= 32'b00111101100000111011101001101111 ;
        1584: q <= 32'b10111101010111010100011001000010 ;
        1585: q <= 32'b00111100101111001111100110110001 ;
        1586: q <= 32'b00111100111110010010010010000010 ;
        1587: q <= 32'b10111101001010110110000010110100 ;
        1588: q <= 32'b10111101100001000101100001011110 ;
        1589: q <= 32'b00111100001001000111110110001111 ;
        1590: q <= 32'b10111101000010001010111101000000 ;
        1591: q <= 32'b10111100001010000100100110001001 ;
        1592: q <= 32'b00111100011000110010000000111101 ;
        1593: q <= 32'b00111101010011110110101111101011 ;
        1594: q <= 32'b10111101100101010110101000000001 ;
        1595: q <= 32'b10111011000011111000001000100110 ;
        1596: q <= 32'b00111100100100110111011101111000 ;
        1597: q <= 32'b10111101110001000111000110110110 ;
        1598: q <= 32'b00111101010010011001001011111010 ;
        1599: q <= 32'b10111101101011000011110100010010 ;
        1600: q <= 32'b10111101010111000111011001010100 ;
        1601: q <= 32'b10111101010000000111011110011101 ;
        1602: q <= 32'b10111101010111111101101111001001 ;
        1603: q <= 32'b00111100101110001011000001011010 ;
        1604: q <= 32'b00111110000101100010011000100110 ;
        1605: q <= 32'b00111101100111011000001110010100 ;
        1606: q <= 32'b10111100001101100111100110000000 ;
        1607: q <= 32'b10111101010000111110110100110100 ;
        1608: q <= 32'b10111110001001110111010111110001 ;
        1609: q <= 32'b00111101011001011101001010100110 ;
        1610: q <= 32'b00111101111000111100000100001100 ;
        1611: q <= 32'b10111011001000110101101001100011 ;
        1612: q <= 32'b10111100010000011000100011011010 ;
        1613: q <= 32'b00111101000011101110101011110001 ;
        1614: q <= 32'b00111100101001111101001001001010 ;
        1615: q <= 32'b10111110000101011011101100010110 ;
        1616: q <= 32'b00111101110000001101011001110011 ;
        1617: q <= 32'b00111110001110111110010010111010 ;
        1618: q <= 32'b00111101110110001000110000001110 ;
        1619: q <= 32'b10111101101100010100101100010110 ;
        1620: q <= 32'b10111101110000110110101011010000 ;
        1621: q <= 32'b10111101101011100011110111010100 ;
        1622: q <= 32'b00111100001111100001101010111000 ;
        1623: q <= 32'b10111100101001111000101110111000 ;
        1624: q <= 32'b10111011100101010000011011111011 ;
        1625: q <= 32'b00111101100011110100101001100011 ;
        1626: q <= 32'b00111011110101000101010001000000 ;
        1627: q <= 32'b10111101001101011111101100101000 ;
        1628: q <= 32'b10111101101110101001001001011011 ;
        1629: q <= 32'b00111100110101110010101010111011 ;
        1630: q <= 32'b00111101100101011011101111011101 ;
        1631: q <= 32'b00111101111101000010111000000100 ;
        1632: q <= 32'b00111101000110001101010001000011 ;
        1633: q <= 32'b00111101110110101110110111001001 ;
        1634: q <= 32'b00111101101011000010000001001011 ;
        1635: q <= 32'b00111110000001111011001000100101 ;
        1636: q <= 32'b10111100100000011001011001011011 ;
        1637: q <= 32'b10111100110100100010010001100100 ;
        1638: q <= 32'b00111110000000011010010100011111 ;
        1639: q <= 32'b10111101011110111111110111110010 ;
        1640: q <= 32'b00000000000000000000000000000000 ;
        1641: q <= 32'b00000000000000000000000000000000 ;
        1642: q <= 32'b00000000000000000000000000000000 ;
        1643: q <= 32'b00000000000000000000000000000000 ;
        1644: q <= 32'b00000000000000000000000000000000 ;
        1645: q <= 32'b00000000000000000000000000000000 ;
        1646: q <= 32'b00000000000000000000000000000000 ;
        1647: q <= 32'b00000000000000000000000000000000 ;
        1648: q <= 32'b00000000000000000000000000000000 ;
        1649: q <= 32'b00000000000000000000000000000000 ;
        1650: q <= 32'b00000000000000000000000000000000 ;
        1651: q <= 32'b00000000000000000000000000000000 ;
        1652: q <= 32'b00000000000000000000000000000000 ;
        1653: q <= 32'b00000000000000000000000000000000 ;
        1654: q <= 32'b00000000000000000000000000000000 ;
        1655: q <= 32'b00000000000000000000000000000000 ;
        1656: q <= 32'b00000000000000000000000000000000 ;
        1657: q <= 32'b00000000000000000000000000000000 ;
        1658: q <= 32'b00000000000000000000000000000000 ;
        1659: q <= 32'b00000000000000000000000000000000 ;
        1660: q <= 32'b00000000000000000000000000000000 ;
        1661: q <= 32'b00000000000000000000000000000000 ;
        1662: q <= 32'b00000000000000000000000000000000 ;
        1663: q <= 32'b00000000000000000000000000000000 ;
        1664: q <= 32'b00111101001000010000010001110100 ;
        1665: q <= 32'b00111101001000000100111100100100 ;
        1666: q <= 32'b10111101011010100110110110010101 ;
        1667: q <= 32'b00111100110001000101001000011111 ;
        1668: q <= 32'b00111101001110101000010010101101 ;
        1669: q <= 32'b00111100111011001010000110001111 ;
        1670: q <= 32'b00111100110010010001101100000111 ;
        1671: q <= 32'b10111100101000011000010101000001 ;
        1672: q <= 32'b10111101010111101100110011101000 ;
        1673: q <= 32'b10111011101000111001011010001011 ;
        1674: q <= 32'b00111101010000001111110010111111 ;
        1675: q <= 32'b00111101101100100111010110101011 ;
        1676: q <= 32'b10111101101001101010000100101110 ;
        1677: q <= 32'b10111101100110001001000011111000 ;
        1678: q <= 32'b00111110000101111010100001001111 ;
        1679: q <= 32'b10111101100010111101100100000100 ;
        1680: q <= 32'b10111101101011011100101000000101 ;
        1681: q <= 32'b00111101010011010010011110011100 ;
        1682: q <= 32'b00111100001100000110000100101111 ;
        1683: q <= 32'b10111101101010100011110101011011 ;
        1684: q <= 32'b10111101110001111000011011101111 ;
        1685: q <= 32'b00111101001111111101100110010000 ;
        1686: q <= 32'b00111100111111110000001101101111 ;
        1687: q <= 32'b00111110000011111100010011011111 ;
        1688: q <= 32'b00111010010101001101101001101111 ;
        1689: q <= 32'b00111100110011010100100000000100 ;
        1690: q <= 32'b10111101110010000000010010100000 ;
        1691: q <= 32'b00111101010110000100000100000000 ;
        1692: q <= 32'b00111100110110011000000010001100 ;
        1693: q <= 32'b10111101111100001001011010110001 ;
        1694: q <= 32'b00111100100110001011100000000001 ;
        1695: q <= 32'b00111101011011010110111010110001 ;
        1696: q <= 32'b00111100010111011001110010011101 ;
        1697: q <= 32'b10111100100100001011101010001001 ;
        1698: q <= 32'b10111101000010011001101100101110 ;
        1699: q <= 32'b00111100111001001001101101111101 ;
        1700: q <= 32'b10111101010011111010001010000101 ;
        1701: q <= 32'b10111100110011001110110101101111 ;
        1702: q <= 32'b00111101101101100101101111001010 ;
        1703: q <= 32'b10111101100110000010101101010100 ;
        1704: q <= 32'b00111101100100100000110010000100 ;
        1705: q <= 32'b00111101011011111111001110110011 ;
        1706: q <= 32'b00111100110110011001100001100100 ;
        1707: q <= 32'b10111101100001010000101100011001 ;
        1708: q <= 32'b00111101110100101110111001001010 ;
        1709: q <= 32'b10111100110100100101000000001100 ;
        1710: q <= 32'b00111101001000010011011111111011 ;
        1711: q <= 32'b00111101110111010111100101001110 ;
        1712: q <= 32'b10111101011100000111000000000010 ;
        1713: q <= 32'b00111101100011011010000110110101 ;
        1714: q <= 32'b10111100000111011000100001001111 ;
        1715: q <= 32'b10111011010011110010101110011001 ;
        1716: q <= 32'b10111110001000110011010110101110 ;
        1717: q <= 32'b00111101011110101110001001000110 ;
        1718: q <= 32'b10111101111001000101010100000111 ;
        1719: q <= 32'b10111101110100010010100110100001 ;
        1720: q <= 32'b10111101101101110101010010010101 ;
        1721: q <= 32'b00111101100101101100011001011000 ;
        1722: q <= 32'b00111101100000011010010000100111 ;
        1723: q <= 32'b10111100011010001110010010100011 ;
        1724: q <= 32'b00111101001101010111101111110111 ;
        1725: q <= 32'b00111101011110101011110001101011 ;
        1726: q <= 32'b10111011111001011110101000111110 ;
        1727: q <= 32'b10111101010100110110001000100011 ;
        1728: q <= 32'b10111100101110100100111011111100 ;
        1729: q <= 32'b00111011111101101011010010111000 ;
        1730: q <= 32'b00111001100011110001000000100110 ;
        1731: q <= 32'b00111101111000001001010001001110 ;
        1732: q <= 32'b10111100110111101011110000000110 ;
        1733: q <= 32'b10111101110001011101010110111101 ;
        1734: q <= 32'b00111101100111000100100011010111 ;
        1735: q <= 32'b00111100101000110100100000001000 ;
        1736: q <= 32'b10111100100010110110111001000011 ;
        1737: q <= 32'b00111101110111000110011011000011 ;
        1738: q <= 32'b10111100011101100010110111000101 ;
        1739: q <= 32'b00111101000110110111111001000011 ;
        1740: q <= 32'b00111101000101011011101100111110 ;
        1741: q <= 32'b00111101001111011111000100101110 ;
        1742: q <= 32'b10111101010100100110101101101000 ;
        1743: q <= 32'b00111101010101000100010111001001 ;
        1744: q <= 32'b10111101011110110111011111010001 ;
        1745: q <= 32'b00111011010000100101101000101011 ;
        1746: q <= 32'b00111101000101101010010101011011 ;
        1747: q <= 32'b10111100100100110000010100110011 ;
        1748: q <= 32'b10111101001110011110010110000110 ;
        1749: q <= 32'b10111100110011100100110111101110 ;
        1750: q <= 32'b10111101010101000111010110101000 ;
        1751: q <= 32'b10111101010000110010111101100011 ;
        1752: q <= 32'b10111100110010101100001001000100 ;
        1753: q <= 32'b10111101000110000000001010011101 ;
        1754: q <= 32'b00111100011100011111001010010000 ;
        1755: q <= 32'b00111101100001110101100001111011 ;
        1756: q <= 32'b00111011011001101110001101111111 ;
        1757: q <= 32'b00111101111011100010001010100010 ;
        1758: q <= 32'b00111101101100110110000101000001 ;
        1759: q <= 32'b00111100011111010010111001101100 ;
        1760: q <= 32'b10111100010010000010010000100010 ;
        1761: q <= 32'b00111100101100101001111100000001 ;
        1762: q <= 32'b10111100010011011000011110100111 ;
        1763: q <= 32'b00111101001101011110110011101010 ;
        1764: q <= 32'b10111101010111100100000010001001 ;
        1765: q <= 32'b10111101101110110001101110001101 ;
        1766: q <= 32'b00111101011101111101001010110000 ;
        1767: q <= 32'b10111101110101011110101010111000 ;
        1768: q <= 32'b00000000000000000000000000000000 ;
        1769: q <= 32'b00000000000000000000000000000000 ;
        1770: q <= 32'b00000000000000000000000000000000 ;
        1771: q <= 32'b00000000000000000000000000000000 ;
        1772: q <= 32'b00000000000000000000000000000000 ;
        1773: q <= 32'b00000000000000000000000000000000 ;
        1774: q <= 32'b00000000000000000000000000000000 ;
        1775: q <= 32'b00000000000000000000000000000000 ;
        1776: q <= 32'b00000000000000000000000000000000 ;
        1777: q <= 32'b00000000000000000000000000000000 ;
        1778: q <= 32'b00000000000000000000000000000000 ;
        1779: q <= 32'b00000000000000000000000000000000 ;
        1780: q <= 32'b00000000000000000000000000000000 ;
        1781: q <= 32'b00000000000000000000000000000000 ;
        1782: q <= 32'b00000000000000000000000000000000 ;
        1783: q <= 32'b00000000000000000000000000000000 ;
        1784: q <= 32'b00000000000000000000000000000000 ;
        1785: q <= 32'b00000000000000000000000000000000 ;
        1786: q <= 32'b00000000000000000000000000000000 ;
        1787: q <= 32'b00000000000000000000000000000000 ;
        1788: q <= 32'b00000000000000000000000000000000 ;
        1789: q <= 32'b00000000000000000000000000000000 ;
        1790: q <= 32'b00000000000000000000000000000000 ;
        1791: q <= 32'b00000000000000000000000000000000 ;
        1792: q <= 32'b10111100000011100001100001110100 ;
        1793: q <= 32'b10111110001011100010010100010100 ;
        1794: q <= 32'b10111101010110111011110111011000 ;
        1795: q <= 32'b00111101001100011100111010000101 ;
        1796: q <= 32'b00111101000101001010010111010001 ;
        1797: q <= 32'b00111101011101110110101110110011 ;
        1798: q <= 32'b00111101111010000100010110000111 ;
        1799: q <= 32'b00111100111101011001110110100010 ;
        1800: q <= 32'b10111101001111100111001011010101 ;
        1801: q <= 32'b00111101010100110010110110010001 ;
        1802: q <= 32'b00111100001001111010111110101100 ;
        1803: q <= 32'b00111101001110110100110011101000 ;
        1804: q <= 32'b10111101100111111011100101001110 ;
        1805: q <= 32'b00111101100101000001000110010010 ;
        1806: q <= 32'b10111101100010110001001010010011 ;
        1807: q <= 32'b00111101100111100100110110111101 ;
        1808: q <= 32'b10111101001100011100101101001001 ;
        1809: q <= 32'b00111101100110111110001110111100 ;
        1810: q <= 32'b10111101111001100010010111111100 ;
        1811: q <= 32'b00111101001100111011101111101011 ;
        1812: q <= 32'b00111101101000110100111000110011 ;
        1813: q <= 32'b10111101010111001100011011101100 ;
        1814: q <= 32'b10111101100000111111111101110110 ;
        1815: q <= 32'b00111101011000001101111110110011 ;
        1816: q <= 32'b10111101100111111111110111001110 ;
        1817: q <= 32'b10111101010001110100011111011111 ;
        1818: q <= 32'b00111011011110000010010111101101 ;
        1819: q <= 32'b10111101101000010001011010011111 ;
        1820: q <= 32'b00111100010000111010001100001011 ;
        1821: q <= 32'b00111101111101111011010001011101 ;
        1822: q <= 32'b10111101010100010101110011101010 ;
        1823: q <= 32'b10111101010110100010110110000000 ;
        1824: q <= 32'b00111101101001001100011111001000 ;
        1825: q <= 32'b00111101001000110001110010000000 ;
        1826: q <= 32'b00111100100000000111010000101101 ;
        1827: q <= 32'b00111101001110110011001111010101 ;
        1828: q <= 32'b00111101001111000010111111001111 ;
        1829: q <= 32'b00111100001100100000100101101001 ;
        1830: q <= 32'b10111101010100100000100010001001 ;
        1831: q <= 32'b10111101110000110110000110000101 ;
        1832: q <= 32'b10111100100011101000100111011010 ;
        1833: q <= 32'b00111100111000100111111011111011 ;
        1834: q <= 32'b00111101100010000110101110010010 ;
        1835: q <= 32'b00111101000100100111110111111111 ;
        1836: q <= 32'b00111100111101111010000000110101 ;
        1837: q <= 32'b10111101010010111101100000000010 ;
        1838: q <= 32'b10111101100111111011011010100000 ;
        1839: q <= 32'b00111100001110000011111010101110 ;
        1840: q <= 32'b10111101100111000111111110000000 ;
        1841: q <= 32'b00111001101111100101000011101110 ;
        1842: q <= 32'b10111100100100000110110111010110 ;
        1843: q <= 32'b00111101010011001001011011001101 ;
        1844: q <= 32'b00111100100011100110110101001101 ;
        1845: q <= 32'b10111101100010101100001001101110 ;
        1846: q <= 32'b10111101111011010111010000001011 ;
        1847: q <= 32'b00111101111100001110010010001111 ;
        1848: q <= 32'b00111100010101010110110011000100 ;
        1849: q <= 32'b10111101111100001001111011000111 ;
        1850: q <= 32'b00111101000000110001000001011100 ;
        1851: q <= 32'b00111100101010011001001011000000 ;
        1852: q <= 32'b00111011100000101110101001100110 ;
        1853: q <= 32'b00111101000001110111101000100110 ;
        1854: q <= 32'b10111101001011110011111000011011 ;
        1855: q <= 32'b00111011100001100101100000111011 ;
        1856: q <= 32'b10111101010001000011100110100101 ;
        1857: q <= 32'b10111101101111001001010010000101 ;
        1858: q <= 32'b10111101101100110001101100110100 ;
        1859: q <= 32'b10111100110110000110010010011010 ;
        1860: q <= 32'b10111100011111010110100011001100 ;
        1861: q <= 32'b00111110001011001111011101001110 ;
        1862: q <= 32'b00111100101011100111100100000101 ;
        1863: q <= 32'b10111110001101001111011010101011 ;
        1864: q <= 32'b10111101010110110110101100010010 ;
        1865: q <= 32'b10111100010101110100101000110001 ;
        1866: q <= 32'b10111110001010001001011010101111 ;
        1867: q <= 32'b00111101110001001111000111111111 ;
        1868: q <= 32'b00111100111001110000100010111101 ;
        1869: q <= 32'b00111101101010100010010001011011 ;
        1870: q <= 32'b10111010100000101100100110011001 ;
        1871: q <= 32'b10111101111101001111111111011101 ;
        1872: q <= 32'b10111101000101001101100000100101 ;
        1873: q <= 32'b10111101100110011010000110001101 ;
        1874: q <= 32'b00111101010000011110001101010000 ;
        1875: q <= 32'b10111110000011111010111110110111 ;
        1876: q <= 32'b10111101111100101001010111001010 ;
        1877: q <= 32'b10111101011001101010011110011001 ;
        1878: q <= 32'b00111100110111010101011100110000 ;
        1879: q <= 32'b10111101011000110001100001011100 ;
        1880: q <= 32'b10111101100111010101010000011111 ;
        1881: q <= 32'b00111101101011011110101110101111 ;
        1882: q <= 32'b10111100011010100101011111110011 ;
        1883: q <= 32'b10111110001101101110111110011011 ;
        1884: q <= 32'b10111101101010011110111110010011 ;
        1885: q <= 32'b00111101011001100101110100000110 ;
        1886: q <= 32'b10111101100000000101101000111001 ;
        1887: q <= 32'b10111101011111001010110100111010 ;
        1888: q <= 32'b00111101001000000010111111011101 ;
        1889: q <= 32'b00111101000110101001011010000110 ;
        1890: q <= 32'b10111100100101011000001000001101 ;
        1891: q <= 32'b10111100110111111101010010101101 ;
        1892: q <= 32'b10111100001100011010100100011110 ;
        1893: q <= 32'b10111101100111110010010001100000 ;
        1894: q <= 32'b00111101000011110001001101000001 ;
        1895: q <= 32'b10111101100001101111101000111000 ;
        1896: q <= 32'b00000000000000000000000000000000 ;
        1897: q <= 32'b00000000000000000000000000000000 ;
        1898: q <= 32'b00000000000000000000000000000000 ;
        1899: q <= 32'b00000000000000000000000000000000 ;
        1900: q <= 32'b00000000000000000000000000000000 ;
        1901: q <= 32'b00000000000000000000000000000000 ;
        1902: q <= 32'b00000000000000000000000000000000 ;
        1903: q <= 32'b00000000000000000000000000000000 ;
        1904: q <= 32'b00000000000000000000000000000000 ;
        1905: q <= 32'b00000000000000000000000000000000 ;
        1906: q <= 32'b00000000000000000000000000000000 ;
        1907: q <= 32'b00000000000000000000000000000000 ;
        1908: q <= 32'b00000000000000000000000000000000 ;
        1909: q <= 32'b00000000000000000000000000000000 ;
        1910: q <= 32'b00000000000000000000000000000000 ;
        1911: q <= 32'b00000000000000000000000000000000 ;
        1912: q <= 32'b00000000000000000000000000000000 ;
        1913: q <= 32'b00000000000000000000000000000000 ;
        1914: q <= 32'b00000000000000000000000000000000 ;
        1915: q <= 32'b00000000000000000000000000000000 ;
        1916: q <= 32'b00000000000000000000000000000000 ;
        1917: q <= 32'b00000000000000000000000000000000 ;
        1918: q <= 32'b00000000000000000000000000000000 ;
        1919: q <= 32'b00000000000000000000000000000000 ;
        1920: q <= 32'b00111100111011011100000010010100 ;
        1921: q <= 32'b10111101101011100001001010010010 ;
        1922: q <= 32'b00111100101011001010010011110000 ;
        1923: q <= 32'b10111100001101101010000001110010 ;
        1924: q <= 32'b00111101100011001111001000101101 ;
        1925: q <= 32'b00111100001010010010101100111010 ;
        1926: q <= 32'b00111011001000100110011011100010 ;
        1927: q <= 32'b10111101101110100000001100011101 ;
        1928: q <= 32'b10111101010101110111101010110101 ;
        1929: q <= 32'b10111101011101111110000100101111 ;
        1930: q <= 32'b10111101100110011000110001110100 ;
        1931: q <= 32'b00111100111100001001011001000100 ;
        1932: q <= 32'b00111100001111011111001111111111 ;
        1933: q <= 32'b10111101100001110110001111110011 ;
        1934: q <= 32'b10111101000100111100111001011111 ;
        1935: q <= 32'b10111101100010000100110110001011 ;
        1936: q <= 32'b00111110000100011010001100000110 ;
        1937: q <= 32'b10111101110010111100110111001001 ;
        1938: q <= 32'b00111100010100000010010011110111 ;
        1939: q <= 32'b00111101110101011001001111100110 ;
        1940: q <= 32'b10111011111100010010001101111000 ;
        1941: q <= 32'b10111100001101010011101001111010 ;
        1942: q <= 32'b10111101101100000111011110101110 ;
        1943: q <= 32'b10111011001000100011110011010001 ;
        1944: q <= 32'b10111101000010111010011010010101 ;
        1945: q <= 32'b10111101100001101111001111101011 ;
        1946: q <= 32'b10111101010011010011111110100011 ;
        1947: q <= 32'b10111110000111111000100111100011 ;
        1948: q <= 32'b10111101110100110110011111010100 ;
        1949: q <= 32'b00111101000101011100100010010001 ;
        1950: q <= 32'b00111100010100011101110111111100 ;
        1951: q <= 32'b00111101010011101001011101000000 ;
        1952: q <= 32'b10111101001000111100010010111110 ;
        1953: q <= 32'b00111100101001000100110000111101 ;
        1954: q <= 32'b10111100110111010111110000011110 ;
        1955: q <= 32'b10111101001010000000110001100110 ;
        1956: q <= 32'b00111100011111100110101000011111 ;
        1957: q <= 32'b00111101001010000010111100011010 ;
        1958: q <= 32'b00111100001010111111011011011010 ;
        1959: q <= 32'b10111101110111001001100010100100 ;
        1960: q <= 32'b00111101000010011010101000001111 ;
        1961: q <= 32'b10111100010011111100110001010010 ;
        1962: q <= 32'b10111101100110101110101000001000 ;
        1963: q <= 32'b10111100100000010100101111110110 ;
        1964: q <= 32'b10111100011011100001010110011101 ;
        1965: q <= 32'b10111101001000110111100111100010 ;
        1966: q <= 32'b10111101000100111101110000100000 ;
        1967: q <= 32'b10111101101011011010111011011100 ;
        1968: q <= 32'b10111101000101100110100000111011 ;
        1969: q <= 32'b10111101000100000000100011101100 ;
        1970: q <= 32'b00111100011000001001111011111001 ;
        1971: q <= 32'b00111101101011001101110100001100 ;
        1972: q <= 32'b10111011000101001011100110010110 ;
        1973: q <= 32'b10111101011000000100111001111101 ;
        1974: q <= 32'b00111101010000010001111111011111 ;
        1975: q <= 32'b00111101101011000011011110010000 ;
        1976: q <= 32'b10111100100110111010101001010110 ;
        1977: q <= 32'b00111100001110000111011101111111 ;
        1978: q <= 32'b00111101111010101100101001010000 ;
        1979: q <= 32'b00111101100000010011010000111111 ;
        1980: q <= 32'b00111100000101111000010010011000 ;
        1981: q <= 32'b10111100111001110100001001101110 ;
        1982: q <= 32'b00111100100101111001101000100010 ;
        1983: q <= 32'b00111101010000111110001000111111 ;
        1984: q <= 32'b00111101101001001011000100000011 ;
        1985: q <= 32'b10111101101100001001010111010001 ;
        1986: q <= 32'b00111101100110011101100100000000 ;
        1987: q <= 32'b00111101101100000001111011111110 ;
        1988: q <= 32'b10111101111010011010001001110100 ;
        1989: q <= 32'b10111101100100000010010111010011 ;
        1990: q <= 32'b10111101101000000000111111001010 ;
        1991: q <= 32'b00111101101001101101010111011110 ;
        1992: q <= 32'b10111011000000101111111011110000 ;
        1993: q <= 32'b10111101000010101100100010111001 ;
        1994: q <= 32'b00111101100001011011001001010101 ;
        1995: q <= 32'b00111101001010000101001110111000 ;
        1996: q <= 32'b10111101101000011000101010100011 ;
        1997: q <= 32'b00111100010011001100000111111111 ;
        1998: q <= 32'b00111101000110000111101100010100 ;
        1999: q <= 32'b10111110000101010111011110110111 ;
        2000: q <= 32'b00111100101011101101111010010000 ;
        2001: q <= 32'b10111101011010010100110100111001 ;
        2002: q <= 32'b00111110000001011101010101100000 ;
        2003: q <= 32'b00111101010001010000110111100001 ;
        2004: q <= 32'b00111101101100010110010100010010 ;
        2005: q <= 32'b10111101100000101111100100000111 ;
        2006: q <= 32'b00111101001010101010010111110110 ;
        2007: q <= 32'b00111101010101101000010111100000 ;
        2008: q <= 32'b00111101000111011111011000000101 ;
        2009: q <= 32'b10111101100000110000101000010010 ;
        2010: q <= 32'b00111101100000001111110000101000 ;
        2011: q <= 32'b00111101001101000110110001111101 ;
        2012: q <= 32'b00111101001100000100111010100010 ;
        2013: q <= 32'b00111101110000100011111011110000 ;
        2014: q <= 32'b10111101100101011110000100110111 ;
        2015: q <= 32'b00111101001001101001111100010110 ;
        2016: q <= 32'b10111101111101001000101000011110 ;
        2017: q <= 32'b10111101011101000010000011011000 ;
        2018: q <= 32'b10111100000110000111100011011111 ;
        2019: q <= 32'b00111100110110101111011111011110 ;
        2020: q <= 32'b10111100100001110000111010111110 ;
        2021: q <= 32'b10111101100011101100010010011010 ;
        2022: q <= 32'b00111101010100111101111100100001 ;
        2023: q <= 32'b00111010111101110101110111010111 ;
        2024: q <= 32'b00000000000000000000000000000000 ;
        2025: q <= 32'b00000000000000000000000000000000 ;
        2026: q <= 32'b00000000000000000000000000000000 ;
        2027: q <= 32'b00000000000000000000000000000000 ;
        2028: q <= 32'b00000000000000000000000000000000 ;
        2029: q <= 32'b00000000000000000000000000000000 ;
        2030: q <= 32'b00000000000000000000000000000000 ;
        2031: q <= 32'b00000000000000000000000000000000 ;
        2032: q <= 32'b00000000000000000000000000000000 ;
        2033: q <= 32'b00000000000000000000000000000000 ;
        2034: q <= 32'b00000000000000000000000000000000 ;
        2035: q <= 32'b00000000000000000000000000000000 ;
        2036: q <= 32'b00000000000000000000000000000000 ;
        2037: q <= 32'b00000000000000000000000000000000 ;
        2038: q <= 32'b00000000000000000000000000000000 ;
        2039: q <= 32'b00000000000000000000000000000000 ;
        2040: q <= 32'b00000000000000000000000000000000 ;
        2041: q <= 32'b00000000000000000000000000000000 ;
        2042: q <= 32'b00000000000000000000000000000000 ;
        2043: q <= 32'b00000000000000000000000000000000 ;
        2044: q <= 32'b00000000000000000000000000000000 ;
        2045: q <= 32'b00000000000000000000000000000000 ;
        2046: q <= 32'b00000000000000000000000000000000 ;
        2047: q <= 32'b00000000000000000000000000000000 ;
        2048: q <= 32'b10111011101001011011101101110000 ;
        2049: q <= 32'b00111101110000110110010111011011 ;
        2050: q <= 32'b00111101010110111001001010111100 ;
        2051: q <= 32'b10111100010101010111111100011110 ;
        2052: q <= 32'b10111101010000111100011000000110 ;
        2053: q <= 32'b10111101101010011111011010001001 ;
        2054: q <= 32'b00111101100010100100111010110110 ;
        2055: q <= 32'b10111101100010111110011111110110 ;
        2056: q <= 32'b10111101001001111111010001000011 ;
        2057: q <= 32'b00111101110010010010111100101100 ;
        2058: q <= 32'b10111100111001111001000000000101 ;
        2059: q <= 32'b10111011110100101100000111100000 ;
        2060: q <= 32'b00111101100110101001010010110100 ;
        2061: q <= 32'b10111110000010101011100111010110 ;
        2062: q <= 32'b10111101110001001011111011011100 ;
        2063: q <= 32'b00111100110001010011000001101011 ;
        2064: q <= 32'b00111100111100001110011110110101 ;
        2065: q <= 32'b00111100000110110100100001101011 ;
        2066: q <= 32'b10111101100100011100100000000111 ;
        2067: q <= 32'b00111101101011101110100111100000 ;
        2068: q <= 32'b00111101100101000100011110110110 ;
        2069: q <= 32'b10111011000100100011101111001111 ;
        2070: q <= 32'b10111110000001110000111001010000 ;
        2071: q <= 32'b10111110000011101101011101010111 ;
        2072: q <= 32'b00111101111110111101010111010000 ;
        2073: q <= 32'b00111101100110011010110100100010 ;
        2074: q <= 32'b00111101101000001010000011111011 ;
        2075: q <= 32'b10111011110111010011001100010001 ;
        2076: q <= 32'b10111101110101001101001111101000 ;
        2077: q <= 32'b00111101001110101000011110011010 ;
        2078: q <= 32'b00111001001001001111001101001000 ;
        2079: q <= 32'b10111100110101100011101111010110 ;
        2080: q <= 32'b00111101110010001001000110000111 ;
        2081: q <= 32'b00111101111011000000110010001110 ;
        2082: q <= 32'b10111101101101001010011100011011 ;
        2083: q <= 32'b00111101101101000100001100000011 ;
        2084: q <= 32'b10111101111010100000101001010110 ;
        2085: q <= 32'b00111100000100111001010100101011 ;
        2086: q <= 32'b10111101101101111010001001110100 ;
        2087: q <= 32'b10111101000001000100100001010000 ;
        2088: q <= 32'b00111101001101001111111110010010 ;
        2089: q <= 32'b10111101111001011011010000101110 ;
        2090: q <= 32'b10111101011001111111001101011110 ;
        2091: q <= 32'b00111110001110101011000100110010 ;
        2092: q <= 32'b10111110000011101001010101001111 ;
        2093: q <= 32'b10111101000001110101000100110001 ;
        2094: q <= 32'b00111101001110111000111111011011 ;
        2095: q <= 32'b10111101100101111001011011101111 ;
        2096: q <= 32'b00111101000000001101110100101001 ;
        2097: q <= 32'b10111101101001010000110100101100 ;
        2098: q <= 32'b10111100110111110011001110011111 ;
        2099: q <= 32'b10111101000010100110101001011010 ;
        2100: q <= 32'b00111101011001011100000111111010 ;
        2101: q <= 32'b00111101100001110100100000001101 ;
        2102: q <= 32'b10111010101111001110111010100000 ;
        2103: q <= 32'b10111101001101111110010101000000 ;
        2104: q <= 32'b00111101001011110101111001001100 ;
        2105: q <= 32'b00111100110110101011001000010110 ;
        2106: q <= 32'b00111101101101011000000110001000 ;
        2107: q <= 32'b00111101101010000100010111111011 ;
        2108: q <= 32'b00111100100101010100011001011101 ;
        2109: q <= 32'b10111011100011101110110011110011 ;
        2110: q <= 32'b00111101101100011111110011100000 ;
        2111: q <= 32'b00111010100000110111111010110000 ;
        2112: q <= 32'b10111100110000110010101101011111 ;
        2113: q <= 32'b00111101011001000001000001001100 ;
        2114: q <= 32'b00111101110001000111000100010110 ;
        2115: q <= 32'b10111101111001101100100001010110 ;
        2116: q <= 32'b00111100111101001000001110110100 ;
        2117: q <= 32'b00111101110100000100101011010000 ;
        2118: q <= 32'b10111011001110101001101111100010 ;
        2119: q <= 32'b00111101000110111000001011010110 ;
        2120: q <= 32'b00111100011100010110000000101101 ;
        2121: q <= 32'b00111101100101001110000011110110 ;
        2122: q <= 32'b10111101000011000101110010000101 ;
        2123: q <= 32'b10111011111110101110100100101111 ;
        2124: q <= 32'b00111101101000001111011001011000 ;
        2125: q <= 32'b00111101111011010010011011101011 ;
        2126: q <= 32'b10111100001101100110100111110001 ;
        2127: q <= 32'b00111110001010101110110110100000 ;
        2128: q <= 32'b10111110011100010010000111100000 ;
        2129: q <= 32'b00111101100001100000111011110111 ;
        2130: q <= 32'b00111101011001000000110011001100 ;
        2131: q <= 32'b00111101110000011100001110111010 ;
        2132: q <= 32'b00111101101011011011110101100000 ;
        2133: q <= 32'b10111101010011100101010010110101 ;
        2134: q <= 32'b10111101010010100011001001111100 ;
        2135: q <= 32'b10111101100001101111110111111111 ;
        2136: q <= 32'b00111101101101100001010101101111 ;
        2137: q <= 32'b00111110001100101111001100100011 ;
        2138: q <= 32'b00111101011111101001000111110000 ;
        2139: q <= 32'b00111110000010000110010011010011 ;
        2140: q <= 32'b00111001110111000001010100101100 ;
        2141: q <= 32'b10111101101011000100100010101010 ;
        2142: q <= 32'b00111010001010000101111100000001 ;
        2143: q <= 32'b00111101001101100011001100011101 ;
        2144: q <= 32'b00111101101010101010010111001010 ;
        2145: q <= 32'b00111101000001110011010110101101 ;
        2146: q <= 32'b10111010111010011010100001100111 ;
        2147: q <= 32'b00111101010011011000111110101010 ;
        2148: q <= 32'b10111101101000101000110111111000 ;
        2149: q <= 32'b00111101100101010111101011010101 ;
        2150: q <= 32'b00111101011011101110111001100010 ;
        2151: q <= 32'b10111100011001100100011001011110 ;
        2152: q <= 32'b00000000000000000000000000000000 ;
        2153: q <= 32'b00000000000000000000000000000000 ;
        2154: q <= 32'b00000000000000000000000000000000 ;
        2155: q <= 32'b00000000000000000000000000000000 ;
        2156: q <= 32'b00000000000000000000000000000000 ;
        2157: q <= 32'b00000000000000000000000000000000 ;
        2158: q <= 32'b00000000000000000000000000000000 ;
        2159: q <= 32'b00000000000000000000000000000000 ;
        2160: q <= 32'b00000000000000000000000000000000 ;
        2161: q <= 32'b00000000000000000000000000000000 ;
        2162: q <= 32'b00000000000000000000000000000000 ;
        2163: q <= 32'b00000000000000000000000000000000 ;
        2164: q <= 32'b00000000000000000000000000000000 ;
        2165: q <= 32'b00000000000000000000000000000000 ;
        2166: q <= 32'b00000000000000000000000000000000 ;
        2167: q <= 32'b00000000000000000000000000000000 ;
        2168: q <= 32'b00000000000000000000000000000000 ;
        2169: q <= 32'b00000000000000000000000000000000 ;
        2170: q <= 32'b00000000000000000000000000000000 ;
        2171: q <= 32'b00000000000000000000000000000000 ;
        2172: q <= 32'b00000000000000000000000000000000 ;
        2173: q <= 32'b00000000000000000000000000000000 ;
        2174: q <= 32'b00000000000000000000000000000000 ;
        2175: q <= 32'b00000000000000000000000000000000 ;
        2176: q <= 32'b10111101100101101011101101010100 ;
        2177: q <= 32'b10111101110000101010001110111110 ;
        2178: q <= 32'b10111101101110001011100010001100 ;
        2179: q <= 32'b00111101110000111100100010010010 ;
        2180: q <= 32'b00111110000001110000001101011011 ;
        2181: q <= 32'b00111000001010010011100111111111 ;
        2182: q <= 32'b10111101010011011000011111100101 ;
        2183: q <= 32'b10111100011100110010011101101110 ;
        2184: q <= 32'b10111110000110111011110100100100 ;
        2185: q <= 32'b00111110000000001101000011100111 ;
        2186: q <= 32'b00111101001010110101100100100010 ;
        2187: q <= 32'b10111101100001110111011111110010 ;
        2188: q <= 32'b00111101100111010100100001111010 ;
        2189: q <= 32'b00111100011111000101101100001010 ;
        2190: q <= 32'b10111011001101010001000010001100 ;
        2191: q <= 32'b10111110100010101101101011101011 ;
        2192: q <= 32'b10111101011100001001010001111011 ;
        2193: q <= 32'b00111101100001110010100100110001 ;
        2194: q <= 32'b00111011111010111001100001111110 ;
        2195: q <= 32'b00111101010001001110001010110111 ;
        2196: q <= 32'b00111101010011101100101001000010 ;
        2197: q <= 32'b00111101111101110010110101101001 ;
        2198: q <= 32'b00111101110110011010001001111000 ;
        2199: q <= 32'b10111100100001001001110101100000 ;
        2200: q <= 32'b10111101001110000001101111110100 ;
        2201: q <= 32'b00111101100000110100001101000100 ;
        2202: q <= 32'b10111100110111110010001111110111 ;
        2203: q <= 32'b00111101010000011100001010110011 ;
        2204: q <= 32'b10111101100010010010110100101001 ;
        2205: q <= 32'b00111101111110111101001011000000 ;
        2206: q <= 32'b00111100000100010111001101101001 ;
        2207: q <= 32'b10111101001011101001101000111001 ;
        2208: q <= 32'b10111101100110100101001011010100 ;
        2209: q <= 32'b10111101100100100000010101111001 ;
        2210: q <= 32'b10111100001010001010101100000101 ;
        2211: q <= 32'b00111101111100100010001000101000 ;
        2212: q <= 32'b10111101001011011110011000000100 ;
        2213: q <= 32'b00111100000100000100011000100000 ;
        2214: q <= 32'b10111101110001011000110101101011 ;
        2215: q <= 32'b00111110001001010011100011011101 ;
        2216: q <= 32'b10111101110001100110110011010010 ;
        2217: q <= 32'b10111101011001101100110001101110 ;
        2218: q <= 32'b00111101101010111101000110001111 ;
        2219: q <= 32'b10111100100100101001011111100100 ;
        2220: q <= 32'b10111101010001011001000100001001 ;
        2221: q <= 32'b00111110001101100101111111010000 ;
        2222: q <= 32'b00111100110000001111100101110011 ;
        2223: q <= 32'b00111101011110111110011100101010 ;
        2224: q <= 32'b10111101100111000101100001111110 ;
        2225: q <= 32'b00111101000001111111101110001011 ;
        2226: q <= 32'b10111101100101100101000010010110 ;
        2227: q <= 32'b00111101001000001001101111100111 ;
        2228: q <= 32'b00111101011011101001110010011000 ;
        2229: q <= 32'b00111011100110100001010110000110 ;
        2230: q <= 32'b10111101100011100011011001101111 ;
        2231: q <= 32'b00111101001100101000101110111110 ;
        2232: q <= 32'b00111110000110001010111111000000 ;
        2233: q <= 32'b10111110001101110111100101011111 ;
        2234: q <= 32'b10111101000101110101111100110010 ;
        2235: q <= 32'b00111100110011100100100011000110 ;
        2236: q <= 32'b10111100110111100000011001010011 ;
        2237: q <= 32'b00111101001110001000001101000111 ;
        2238: q <= 32'b10111101001111010101110010000110 ;
        2239: q <= 32'b10111101110011011010010111000011 ;
        2240: q <= 32'b10111101110110101100111000100101 ;
        2241: q <= 32'b00111101011101100001100010001000 ;
        2242: q <= 32'b10111101101010111101111000111111 ;
        2243: q <= 32'b00111011001110101001111100010101 ;
        2244: q <= 32'b10111101011011001000100101111011 ;
        2245: q <= 32'b00111101111100000011001101011000 ;
        2246: q <= 32'b00111100110110110010111001100100 ;
        2247: q <= 32'b00111101110011001000000101111100 ;
        2248: q <= 32'b00111101001111011010000010101111 ;
        2249: q <= 32'b00111110000100001101000100111000 ;
        2250: q <= 32'b10111101100001110011011011000111 ;
        2251: q <= 32'b10111101010000010010010110010011 ;
        2252: q <= 32'b00111101101011000111011111110000 ;
        2253: q <= 32'b10111101101001000101100100011101 ;
        2254: q <= 32'b00111101110101100101011010010111 ;
        2255: q <= 32'b10111101111000011110000100000111 ;
        2256: q <= 32'b10111110000001101000111010101001 ;
        2257: q <= 32'b00111110000100111110001001010111 ;
        2258: q <= 32'b00111101110010111010010111010100 ;
        2259: q <= 32'b10111110000100010000011000110100 ;
        2260: q <= 32'b00111100001100111111101001011011 ;
        2261: q <= 32'b00111101011010100100001101011101 ;
        2262: q <= 32'b10111100000100000000110000110010 ;
        2263: q <= 32'b10111101010100000011110000111100 ;
        2264: q <= 32'b00111101001011111101111001101100 ;
        2265: q <= 32'b00111101001011000000100000100010 ;
        2266: q <= 32'b00111101100100111101110111011010 ;
        2267: q <= 32'b00111011110100101001111010001010 ;
        2268: q <= 32'b10111100010011011101010110111111 ;
        2269: q <= 32'b00111101001000111001100100101100 ;
        2270: q <= 32'b00111100111101011101110001100000 ;
        2271: q <= 32'b00111110001110100011010101111011 ;
        2272: q <= 32'b00111101000100010011101000010111 ;
        2273: q <= 32'b10111100111100011100010100111010 ;
        2274: q <= 32'b00111110010001000010000111010111 ;
        2275: q <= 32'b00111101110100010011011011000000 ;
        2276: q <= 32'b00111101010110001011000110100000 ;
        2277: q <= 32'b00111101111100101110000010011011 ;
        2278: q <= 32'b00111101110000101000011000000101 ;
        2279: q <= 32'b10111101101011101111000001001001 ;
        2280: q <= 32'b00000000000000000000000000000000 ;
        2281: q <= 32'b00000000000000000000000000000000 ;
        2282: q <= 32'b00000000000000000000000000000000 ;
        2283: q <= 32'b00000000000000000000000000000000 ;
        2284: q <= 32'b00000000000000000000000000000000 ;
        2285: q <= 32'b00000000000000000000000000000000 ;
        2286: q <= 32'b00000000000000000000000000000000 ;
        2287: q <= 32'b00000000000000000000000000000000 ;
        2288: q <= 32'b00000000000000000000000000000000 ;
        2289: q <= 32'b00000000000000000000000000000000 ;
        2290: q <= 32'b00000000000000000000000000000000 ;
        2291: q <= 32'b00000000000000000000000000000000 ;
        2292: q <= 32'b00000000000000000000000000000000 ;
        2293: q <= 32'b00000000000000000000000000000000 ;
        2294: q <= 32'b00000000000000000000000000000000 ;
        2295: q <= 32'b00000000000000000000000000000000 ;
        2296: q <= 32'b00000000000000000000000000000000 ;
        2297: q <= 32'b00000000000000000000000000000000 ;
        2298: q <= 32'b00000000000000000000000000000000 ;
        2299: q <= 32'b00000000000000000000000000000000 ;
        2300: q <= 32'b00000000000000000000000000000000 ;
        2301: q <= 32'b00000000000000000000000000000000 ;
        2302: q <= 32'b00000000000000000000000000000000 ;
        2303: q <= 32'b00000000000000000000000000000000 ;
        2304: q <= 32'b10111110000101011001010111001100 ;
        2305: q <= 32'b10111101101001001010010010011011 ;
        2306: q <= 32'b10111101101011100001101011001111 ;
        2307: q <= 32'b10111101101110111101000101101110 ;
        2308: q <= 32'b00111100001111011011011000011110 ;
        2309: q <= 32'b00111101011100110110111100110101 ;
        2310: q <= 32'b10111011101111111110100100000001 ;
        2311: q <= 32'b00111101001110011111101010011101 ;
        2312: q <= 32'b10111101011000110100011001110011 ;
        2313: q <= 32'b10111101101011001001111001011001 ;
        2314: q <= 32'b10111100110100110010111010000111 ;
        2315: q <= 32'b10111101110000010111100111101111 ;
        2316: q <= 32'b10111101101011111000001111010100 ;
        2317: q <= 32'b10111101011011110100101100001101 ;
        2318: q <= 32'b10111101011100101001010101001101 ;
        2319: q <= 32'b10111101001110011010111010010111 ;
        2320: q <= 32'b10111101000100110111011000101000 ;
        2321: q <= 32'b10111101000100110100110101110101 ;
        2322: q <= 32'b00111100100010000010101110011010 ;
        2323: q <= 32'b10111100010110111000111101110111 ;
        2324: q <= 32'b00111101001000011111100001111101 ;
        2325: q <= 32'b10111100110110111101000000101000 ;
        2326: q <= 32'b10111101001001010000110110110010 ;
        2327: q <= 32'b00111101100011100000110011100010 ;
        2328: q <= 32'b00111100100011110111001110000111 ;
        2329: q <= 32'b00111101101011001110011101101111 ;
        2330: q <= 32'b00111100100111011011000101011101 ;
        2331: q <= 32'b00111101100011110100101001001000 ;
        2332: q <= 32'b00111100111110110100001000000011 ;
        2333: q <= 32'b00111101011011001000110101010001 ;
        2334: q <= 32'b10111101011011000000100000011111 ;
        2335: q <= 32'b10111101010110101101110000010000 ;
        2336: q <= 32'b10111011111001001101110010000000 ;
        2337: q <= 32'b10111101110010010110111000111100 ;
        2338: q <= 32'b00111001111101110100000011011001 ;
        2339: q <= 32'b10111101010000011111100000001010 ;
        2340: q <= 32'b10111101001101100000111010000110 ;
        2341: q <= 32'b10111101011001000111110110010000 ;
        2342: q <= 32'b00111101110110101010010111101011 ;
        2343: q <= 32'b00111101101110101000111000100100 ;
        2344: q <= 32'b00111100011100110101111011110011 ;
        2345: q <= 32'b00111101100000001100001001000011 ;
        2346: q <= 32'b00111101010101100001100111000110 ;
        2347: q <= 32'b00111101010110011111001001100011 ;
        2348: q <= 32'b00111101100100111100010010100011 ;
        2349: q <= 32'b10111101101011111011010011111000 ;
        2350: q <= 32'b10111101110001001001100111101010 ;
        2351: q <= 32'b10111100100000111001100111111010 ;
        2352: q <= 32'b00111101100110001001010000000011 ;
        2353: q <= 32'b00111100111111110000101101010110 ;
        2354: q <= 32'b10111101001110000100100100101101 ;
        2355: q <= 32'b00111101100111110000001100100101 ;
        2356: q <= 32'b10111101110011100111001110010100 ;
        2357: q <= 32'b10111101010100011000000010010111 ;
        2358: q <= 32'b10111100101100110011100110001011 ;
        2359: q <= 32'b00111101011000101011010100111110 ;
        2360: q <= 32'b00111101100000111010001110101000 ;
        2361: q <= 32'b00111100010100101110010001011011 ;
        2362: q <= 32'b00111100101111111101011101010100 ;
        2363: q <= 32'b00111101100010000011000001100100 ;
        2364: q <= 32'b10111101110100001100001010011111 ;
        2365: q <= 32'b10111101100110110000101101000001 ;
        2366: q <= 32'b00111011100001001011100000110010 ;
        2367: q <= 32'b10111101010010110111011100101001 ;
        2368: q <= 32'b10111101011000010101011100001101 ;
        2369: q <= 32'b10111100110011100010110011001011 ;
        2370: q <= 32'b00111100100100001000100001001111 ;
        2371: q <= 32'b00111100001100100011010110100001 ;
        2372: q <= 32'b00111101101011011110011010000101 ;
        2373: q <= 32'b00111101100111110001101101101011 ;
        2374: q <= 32'b00111101101011011011010100111011 ;
        2375: q <= 32'b00111101001100001000011111000110 ;
        2376: q <= 32'b10111100100001010111111010100011 ;
        2377: q <= 32'b00111101011110000100000110010000 ;
        2378: q <= 32'b10111101010000111001100001000100 ;
        2379: q <= 32'b10111101000111010100011101101001 ;
        2380: q <= 32'b10111101101001000011110001101111 ;
        2381: q <= 32'b00111101100110000011110110101010 ;
        2382: q <= 32'b10111100001101011010100001110000 ;
        2383: q <= 32'b00111101100010001001011101101101 ;
        2384: q <= 32'b10111101011110111000010101010101 ;
        2385: q <= 32'b00111100100000111101000001000010 ;
        2386: q <= 32'b00111100100000110011111101011001 ;
        2387: q <= 32'b10111100100100111010010000101001 ;
        2388: q <= 32'b10111101110000000000100101110111 ;
        2389: q <= 32'b00111101100000011001011010010101 ;
        2390: q <= 32'b00111100101001010111110001011110 ;
        2391: q <= 32'b10111101011001110001100111110110 ;
        2392: q <= 32'b10111101100111111000000001011101 ;
        2393: q <= 32'b10111101000011100011101011110100 ;
        2394: q <= 32'b00111100110000101110111011100100 ;
        2395: q <= 32'b10111101010101010010000011100001 ;
        2396: q <= 32'b00111101100111101110000111001100 ;
        2397: q <= 32'b00111101100011101100011100010100 ;
        2398: q <= 32'b10111101011010100001000000000100 ;
        2399: q <= 32'b00111101011101101001000111011111 ;
        2400: q <= 32'b00111101010110101100100101001100 ;
        2401: q <= 32'b00111101000111000110001110010001 ;
        2402: q <= 32'b00111100000111100000111000000000 ;
        2403: q <= 32'b10111101001011110110101001111111 ;
        2404: q <= 32'b10111100000010101010100111101101 ;
        2405: q <= 32'b10111100011101000111001010011001 ;
        2406: q <= 32'b10111100100011001110110000111111 ;
        2407: q <= 32'b10111101011000111101101001011100 ;
        2408: q <= 32'b00000000000000000000000000000000 ;
        2409: q <= 32'b00000000000000000000000000000000 ;
        2410: q <= 32'b00000000000000000000000000000000 ;
        2411: q <= 32'b00000000000000000000000000000000 ;
        2412: q <= 32'b00000000000000000000000000000000 ;
        2413: q <= 32'b00000000000000000000000000000000 ;
        2414: q <= 32'b00000000000000000000000000000000 ;
        2415: q <= 32'b00000000000000000000000000000000 ;
        2416: q <= 32'b00000000000000000000000000000000 ;
        2417: q <= 32'b00000000000000000000000000000000 ;
        2418: q <= 32'b00000000000000000000000000000000 ;
        2419: q <= 32'b00000000000000000000000000000000 ;
        2420: q <= 32'b00000000000000000000000000000000 ;
        2421: q <= 32'b00000000000000000000000000000000 ;
        2422: q <= 32'b00000000000000000000000000000000 ;
        2423: q <= 32'b00000000000000000000000000000000 ;
        2424: q <= 32'b00000000000000000000000000000000 ;
        2425: q <= 32'b00000000000000000000000000000000 ;
        2426: q <= 32'b00000000000000000000000000000000 ;
        2427: q <= 32'b00000000000000000000000000000000 ;
        2428: q <= 32'b00000000000000000000000000000000 ;
        2429: q <= 32'b00000000000000000000000000000000 ;
        2430: q <= 32'b00000000000000000000000000000000 ;
        2431: q <= 32'b00000000000000000000000000000000 ;
        2432: q <= 32'b00111100100111000000000010111001 ;
        2433: q <= 32'b00111101011011001101001101111001 ;
        2434: q <= 32'b00111101001111100001000100100001 ;
        2435: q <= 32'b00111100010100001111011101001010 ;
        2436: q <= 32'b10111101110001110010001111010110 ;
        2437: q <= 32'b10111100011000110010110101000100 ;
        2438: q <= 32'b00111101000111111001001110001110 ;
        2439: q <= 32'b10111101100101110101011000110011 ;
        2440: q <= 32'b00111100100111001010001111001010 ;
        2441: q <= 32'b00111100000100011110000010101101 ;
        2442: q <= 32'b10111100100000110001000110011000 ;
        2443: q <= 32'b10111101010110100101100101110000 ;
        2444: q <= 32'b10111100100101111100010101111111 ;
        2445: q <= 32'b00111011001111010010001110111110 ;
        2446: q <= 32'b10111101001110100011001001101111 ;
        2447: q <= 32'b00111101100110001101000100111010 ;
        2448: q <= 32'b10111101010110101010100100010100 ;
        2449: q <= 32'b10111100110010000000001011101110 ;
        2450: q <= 32'b00111110000000001101111101010011 ;
        2451: q <= 32'b10111100011100100100010111111011 ;
        2452: q <= 32'b10111101001100100011010110111100 ;
        2453: q <= 32'b10111101111011000001100110011110 ;
        2454: q <= 32'b10111101110111001100110000001110 ;
        2455: q <= 32'b00111100100010001000011010111101 ;
        2456: q <= 32'b10111101100011010111001101111000 ;
        2457: q <= 32'b10111100111101101110100100000110 ;
        2458: q <= 32'b10111101010010001101100010011111 ;
        2459: q <= 32'b10111101000010001111110001101001 ;
        2460: q <= 32'b00111011110101100101010110101101 ;
        2461: q <= 32'b10111101101110100000010000111110 ;
        2462: q <= 32'b10111101110100111000110101110001 ;
        2463: q <= 32'b00111101000110100000110100101010 ;
        2464: q <= 32'b00111110001010110100100011011100 ;
        2465: q <= 32'b10111101110111110010010100001011 ;
        2466: q <= 32'b00111101010100110101101011011101 ;
        2467: q <= 32'b10111101100001111001101010010101 ;
        2468: q <= 32'b10111101111011001011011000010101 ;
        2469: q <= 32'b00111101000100110101110000011110 ;
        2470: q <= 32'b10111011000101011110100000100001 ;
        2471: q <= 32'b10111101001111111100010101011010 ;
        2472: q <= 32'b00111101001011010001001011100010 ;
        2473: q <= 32'b10111101100100001101110011000110 ;
        2474: q <= 32'b00111101110010000110110010111010 ;
        2475: q <= 32'b00111110000101010001001110100000 ;
        2476: q <= 32'b00111100111110011001110000110101 ;
        2477: q <= 32'b10111101110110110100100100011110 ;
        2478: q <= 32'b00111101001001101001000111100111 ;
        2479: q <= 32'b00111100000111001111000111011001 ;
        2480: q <= 32'b10111101100101100010010010101110 ;
        2481: q <= 32'b00111100001011101001010111000111 ;
        2482: q <= 32'b10111101001101000101000010001000 ;
        2483: q <= 32'b00111101010010011001111110000011 ;
        2484: q <= 32'b00111101111010110111100001101100 ;
        2485: q <= 32'b00111110001001100101111101011000 ;
        2486: q <= 32'b10111100101110111111101110011110 ;
        2487: q <= 32'b00111100110011011010111001101100 ;
        2488: q <= 32'b10111110000101010001000000000101 ;
        2489: q <= 32'b00111101010010111001010110011001 ;
        2490: q <= 32'b00111101111001101000001000011010 ;
        2491: q <= 32'b00111011000010100100001000101111 ;
        2492: q <= 32'b10111101101101111100110011101110 ;
        2493: q <= 32'b10111101101000110000001101011111 ;
        2494: q <= 32'b10111101110011100010001010110000 ;
        2495: q <= 32'b00111101110100011010010110111010 ;
        2496: q <= 32'b00111101001000110011000010010010 ;
        2497: q <= 32'b00111100000010001000111101100011 ;
        2498: q <= 32'b00111110000011101011011000111001 ;
        2499: q <= 32'b10111110010110110010011010011010 ;
        2500: q <= 32'b10111101000001111010001111010001 ;
        2501: q <= 32'b10111101101101110010110000111111 ;
        2502: q <= 32'b00111101001000101011001100010101 ;
        2503: q <= 32'b00111101101100000110000000011111 ;
        2504: q <= 32'b00111100101100101101110010101100 ;
        2505: q <= 32'b10111101001110101110101001100110 ;
        2506: q <= 32'b10111101011110101000100011010101 ;
        2507: q <= 32'b00111100010001001000110000011000 ;
        2508: q <= 32'b10111010011110010001111001101010 ;
        2509: q <= 32'b00111101010110110000010011001011 ;
        2510: q <= 32'b00111100011111011111011100110000 ;
        2511: q <= 32'b10111101010101010111011010110111 ;
        2512: q <= 32'b00111101001110111011011000011100 ;
        2513: q <= 32'b00111100000110110100110011110010 ;
        2514: q <= 32'b10111101001001101101110101000011 ;
        2515: q <= 32'b00111101110000011010100011001111 ;
        2516: q <= 32'b00111101111111100001111010111110 ;
        2517: q <= 32'b10111101100000111001001100000001 ;
        2518: q <= 32'b00111101001010000010001011100110 ;
        2519: q <= 32'b10111100101110001101001000011001 ;
        2520: q <= 32'b00111101011110111001010001100110 ;
        2521: q <= 32'b10111100100111111111110000010101 ;
        2522: q <= 32'b00111101100011010011101001010010 ;
        2523: q <= 32'b10111101101101011101010111111111 ;
        2524: q <= 32'b10111101001000101111000101110011 ;
        2525: q <= 32'b00111011101001100110001000010110 ;
        2526: q <= 32'b10111100110111110001011111111100 ;
        2527: q <= 32'b10111100110000010001010001100010 ;
        2528: q <= 32'b00111100110010011001100110000011 ;
        2529: q <= 32'b00111101010110100101001011101010 ;
        2530: q <= 32'b10111101011000100100011110010010 ;
        2531: q <= 32'b00111100000010010000100000100001 ;
        2532: q <= 32'b00111101010110110110110011000000 ;
        2533: q <= 32'b00111101100010111000000100000010 ;
        2534: q <= 32'b10111100101011110111000101100000 ;
        2535: q <= 32'b00111100100011100001010110000101 ;
        2536: q <= 32'b00000000000000000000000000000000 ;
        2537: q <= 32'b00000000000000000000000000000000 ;
        2538: q <= 32'b00000000000000000000000000000000 ;
        2539: q <= 32'b00000000000000000000000000000000 ;
        2540: q <= 32'b00000000000000000000000000000000 ;
        2541: q <= 32'b00000000000000000000000000000000 ;
        2542: q <= 32'b00000000000000000000000000000000 ;
        2543: q <= 32'b00000000000000000000000000000000 ;
        2544: q <= 32'b00000000000000000000000000000000 ;
        2545: q <= 32'b00000000000000000000000000000000 ;
        2546: q <= 32'b00000000000000000000000000000000 ;
        2547: q <= 32'b00000000000000000000000000000000 ;
        2548: q <= 32'b00000000000000000000000000000000 ;
        2549: q <= 32'b00000000000000000000000000000000 ;
        2550: q <= 32'b00000000000000000000000000000000 ;
        2551: q <= 32'b00000000000000000000000000000000 ;
        2552: q <= 32'b00000000000000000000000000000000 ;
        2553: q <= 32'b00000000000000000000000000000000 ;
        2554: q <= 32'b00000000000000000000000000000000 ;
        2555: q <= 32'b00000000000000000000000000000000 ;
        2556: q <= 32'b00000000000000000000000000000000 ;
        2557: q <= 32'b00000000000000000000000000000000 ;
        2558: q <= 32'b00000000000000000000000000000000 ;
        2559: q <= 32'b00000000000000000000000000000000 ;
        2560: q <= 32'b10111101010011010001000011000110 ;
        2561: q <= 32'b00111110001011110000010101010101 ;
        2562: q <= 32'b00111100101111100101101101101010 ;
        2563: q <= 32'b10111101011111001000001000011101 ;
        2564: q <= 32'b10111101101011110111011001010100 ;
        2565: q <= 32'b00111101100100111110100001101011 ;
        2566: q <= 32'b10111101101001001110110101000001 ;
        2567: q <= 32'b00111101000010111000010100100000 ;
        2568: q <= 32'b00111101100100110010011110000110 ;
        2569: q <= 32'b00111101100000011100001000100100 ;
        2570: q <= 32'b10111101001110100110101010100111 ;
        2571: q <= 32'b10111101011011011100111001110101 ;
        2572: q <= 32'b10111100101101011101011111001111 ;
        2573: q <= 32'b10111101001111111111110100110010 ;
        2574: q <= 32'b10111110000001010100001001101010 ;
        2575: q <= 32'b00111101110001000101010100111101 ;
        2576: q <= 32'b00111100110001000100000001001110 ;
        2577: q <= 32'b10111100011101011100111101000000 ;
        2578: q <= 32'b00111101100001001010100011010010 ;
        2579: q <= 32'b00111101100010111010100110000110 ;
        2580: q <= 32'b00111101110001011110011001010011 ;
        2581: q <= 32'b10111101001101101000110000110010 ;
        2582: q <= 32'b00111101001101100101000101000011 ;
        2583: q <= 32'b10111101101000011010001010001011 ;
        2584: q <= 32'b00111101101011101100100010101100 ;
        2585: q <= 32'b00111101100100101011001011110110 ;
        2586: q <= 32'b00111011010010100011010110001101 ;
        2587: q <= 32'b00111101101010000100000101101101 ;
        2588: q <= 32'b00111101010110101011101110001100 ;
        2589: q <= 32'b00111100101001010000001001101111 ;
        2590: q <= 32'b10111101111001110001101110101010 ;
        2591: q <= 32'b00111100111001000110001011000000 ;
        2592: q <= 32'b00111100111001000011000110011010 ;
        2593: q <= 32'b10111100011011100001010000110101 ;
        2594: q <= 32'b10111101010000111001001100111111 ;
        2595: q <= 32'b10111101100001010000101111000001 ;
        2596: q <= 32'b10111101101110011010011001001000 ;
        2597: q <= 32'b10111100110110100001101010101100 ;
        2598: q <= 32'b00111011001110001000000010011111 ;
        2599: q <= 32'b00111110000011010011101111000010 ;
        2600: q <= 32'b10111110011110001101010010001001 ;
        2601: q <= 32'b10111110000110100100001111100111 ;
        2602: q <= 32'b10111100000011111010011100111010 ;
        2603: q <= 32'b10111101001101101110010111000110 ;
        2604: q <= 32'b10111100110110001010111100110011 ;
        2605: q <= 32'b00111101101010010100111110111101 ;
        2606: q <= 32'b00111011001011100011101101110001 ;
        2607: q <= 32'b10111110000100000111111110001011 ;
        2608: q <= 32'b00111101001000010011001001101000 ;
        2609: q <= 32'b10111101011111001010011000000110 ;
        2610: q <= 32'b00111100110101100000110101101000 ;
        2611: q <= 32'b00111101000000100010101011000011 ;
        2612: q <= 32'b00111101111100110010100000000111 ;
        2613: q <= 32'b10111100001010001110111110101110 ;
        2614: q <= 32'b00111101001001101111001011001010 ;
        2615: q <= 32'b00111011101110110001000110101100 ;
        2616: q <= 32'b10111101110011100010001100001011 ;
        2617: q <= 32'b00111101111110010010110101101101 ;
        2618: q <= 32'b00111101000111110100010110110111 ;
        2619: q <= 32'b10111101110100110111000001101001 ;
        2620: q <= 32'b10111101011100101101100111010011 ;
        2621: q <= 32'b00111100101101010111100101001111 ;
        2622: q <= 32'b10111101100001001101101101001011 ;
        2623: q <= 32'b00111101000100000010011010111101 ;
        2624: q <= 32'b10111101101110111111011010100111 ;
        2625: q <= 32'b00111110000010000100110011001100 ;
        2626: q <= 32'b10111101010011101111100111010000 ;
        2627: q <= 32'b00111101000011011101101011010111 ;
        2628: q <= 32'b10111101100111101001110010011011 ;
        2629: q <= 32'b10111101100110001000011010010101 ;
        2630: q <= 32'b10111101111001100010010100010101 ;
        2631: q <= 32'b00111101100010110100111110001010 ;
        2632: q <= 32'b10111100011101000100111011100111 ;
        2633: q <= 32'b10111101100001110111010011010101 ;
        2634: q <= 32'b10111101100010010100001110110011 ;
        2635: q <= 32'b00111101101001100000101100011001 ;
        2636: q <= 32'b00111101100010110011110000011011 ;
        2637: q <= 32'b00111101010110010111100111001101 ;
        2638: q <= 32'b10111101100000111100110101000101 ;
        2639: q <= 32'b10111101110101011011101000000011 ;
        2640: q <= 32'b10111100100001111101100001011010 ;
        2641: q <= 32'b10111100101101100010000010110011 ;
        2642: q <= 32'b00111101100001111110101010010111 ;
        2643: q <= 32'b00111100100010110100011101011000 ;
        2644: q <= 32'b00111101011101111010111001000111 ;
        2645: q <= 32'b00111101000000111100101101011010 ;
        2646: q <= 32'b10111101001000111010000001010011 ;
        2647: q <= 32'b10111100100111010011111010011010 ;
        2648: q <= 32'b10111100011100000000110111000011 ;
        2649: q <= 32'b10111100100110011010110100000000 ;
        2650: q <= 32'b00111101001011000011011011100010 ;
        2651: q <= 32'b00111100110010001110010001001101 ;
        2652: q <= 32'b10111101011010000110011111111110 ;
        2653: q <= 32'b10111011010001101111110100011110 ;
        2654: q <= 32'b00111101011000101110000100011001 ;
        2655: q <= 32'b10111100110101000110100101010011 ;
        2656: q <= 32'b10111101110001010000111000010010 ;
        2657: q <= 32'b10111011101011001000001100011000 ;
        2658: q <= 32'b00111100001101110110011010011110 ;
        2659: q <= 32'b00111100101011110011110010000000 ;
        2660: q <= 32'b10111101000110101011000100100110 ;
        2661: q <= 32'b00111101000010110111100001110101 ;
        2662: q <= 32'b10111101011010111011001111011010 ;
        2663: q <= 32'b00111101000110100101111111000010 ;
        2664: q <= 32'b00000000000000000000000000000000 ;
        2665: q <= 32'b00000000000000000000000000000000 ;
        2666: q <= 32'b00000000000000000000000000000000 ;
        2667: q <= 32'b00000000000000000000000000000000 ;
        2668: q <= 32'b00000000000000000000000000000000 ;
        2669: q <= 32'b00000000000000000000000000000000 ;
        2670: q <= 32'b00000000000000000000000000000000 ;
        2671: q <= 32'b00000000000000000000000000000000 ;
        2672: q <= 32'b00000000000000000000000000000000 ;
        2673: q <= 32'b00000000000000000000000000000000 ;
        2674: q <= 32'b00000000000000000000000000000000 ;
        2675: q <= 32'b00000000000000000000000000000000 ;
        2676: q <= 32'b00000000000000000000000000000000 ;
        2677: q <= 32'b00000000000000000000000000000000 ;
        2678: q <= 32'b00000000000000000000000000000000 ;
        2679: q <= 32'b00000000000000000000000000000000 ;
        2680: q <= 32'b00000000000000000000000000000000 ;
        2681: q <= 32'b00000000000000000000000000000000 ;
        2682: q <= 32'b00000000000000000000000000000000 ;
        2683: q <= 32'b00000000000000000000000000000000 ;
        2684: q <= 32'b00000000000000000000000000000000 ;
        2685: q <= 32'b00000000000000000000000000000000 ;
        2686: q <= 32'b00000000000000000000000000000000 ;
        2687: q <= 32'b00000000000000000000000000000000 ;
        2688: q <= 32'b10111101010010100101011000110010 ;
        2689: q <= 32'b10111101100011001100111110100000 ;
        2690: q <= 32'b10111010010010010100011011100100 ;
        2691: q <= 32'b10111101110100100010000111001110 ;
        2692: q <= 32'b10111100110111111000100100001110 ;
        2693: q <= 32'b10111101100111001101001101001101 ;
        2694: q <= 32'b00111101101011001011100100100011 ;
        2695: q <= 32'b00111101100110110011100110100111 ;
        2696: q <= 32'b00111100101011001010110110010100 ;
        2697: q <= 32'b10111101000111011111001110011011 ;
        2698: q <= 32'b10111100100110111000011011001110 ;
        2699: q <= 32'b10111100111011110110000110110110 ;
        2700: q <= 32'b10111011000010101010001000010010 ;
        2701: q <= 32'b00111100101000111111011010000011 ;
        2702: q <= 32'b00111101101111010110110000011100 ;
        2703: q <= 32'b10111101010000101000111100110010 ;
        2704: q <= 32'b10111101110101000101111010001010 ;
        2705: q <= 32'b00111100011100010111001101011001 ;
        2706: q <= 32'b10111101010110011101001110010111 ;
        2707: q <= 32'b10111101000010010000110000100111 ;
        2708: q <= 32'b00111101100010101100100101110101 ;
        2709: q <= 32'b10111101011011110101001111100000 ;
        2710: q <= 32'b10111100110010101011110010000100 ;
        2711: q <= 32'b10111101100111101100000110010001 ;
        2712: q <= 32'b00111100110100000101100100011101 ;
        2713: q <= 32'b10111101010111000111011101111100 ;
        2714: q <= 32'b00111101110100011001101111101011 ;
        2715: q <= 32'b00111010101100010111001000010010 ;
        2716: q <= 32'b10111101010010001111011000110110 ;
        2717: q <= 32'b00111101010110000101010010100110 ;
        2718: q <= 32'b10111101011000011101010110101001 ;
        2719: q <= 32'b10111100100010001110011000101000 ;
        2720: q <= 32'b00111101100111000000010101001110 ;
        2721: q <= 32'b00111101100110101101001110010111 ;
        2722: q <= 32'b00111101110001100000100001110001 ;
        2723: q <= 32'b00111011101111001010001010010011 ;
        2724: q <= 32'b10111101111001010001101011011011 ;
        2725: q <= 32'b10111101101000000111100010011000 ;
        2726: q <= 32'b00111101001001100010110001000011 ;
        2727: q <= 32'b00111100000111111010011000010001 ;
        2728: q <= 32'b00111110000011110010001010000110 ;
        2729: q <= 32'b10111011110100010110100110011001 ;
        2730: q <= 32'b00111101001010010000000000100010 ;
        2731: q <= 32'b00111101001110111101111101000011 ;
        2732: q <= 32'b00111011100010100010010010000011 ;
        2733: q <= 32'b00111100111101101001000010000100 ;
        2734: q <= 32'b10111100110000001011010001011100 ;
        2735: q <= 32'b10111101100100000000111001110110 ;
        2736: q <= 32'b10111101101100010110110001010110 ;
        2737: q <= 32'b00111101010110101010001111110110 ;
        2738: q <= 32'b00111101101000010010010011100000 ;
        2739: q <= 32'b10111100101000010110000011001111 ;
        2740: q <= 32'b00111110000001101101010000001101 ;
        2741: q <= 32'b00111101101110000011000011010111 ;
        2742: q <= 32'b10111100110101111100010100001000 ;
        2743: q <= 32'b00111101010001100001000101101100 ;
        2744: q <= 32'b10111101000000001110011000000010 ;
        2745: q <= 32'b10111100111111100111011000110101 ;
        2746: q <= 32'b00111101100101011110000110110100 ;
        2747: q <= 32'b10111100000110010100110100011001 ;
        2748: q <= 32'b00111101000001010101000011010101 ;
        2749: q <= 32'b10111011101111001011011010011110 ;
        2750: q <= 32'b00111010101001001101110010111010 ;
        2751: q <= 32'b00111011110110100001001011010111 ;
        2752: q <= 32'b10111100110110011101111101100101 ;
        2753: q <= 32'b10111101100101011100101111110111 ;
        2754: q <= 32'b10111101100000111001011001001111 ;
        2755: q <= 32'b00111101000100000110011100011000 ;
        2756: q <= 32'b10111011111110001010000001011001 ;
        2757: q <= 32'b00111101100001101010100110101110 ;
        2758: q <= 32'b10111011110110101001100111010111 ;
        2759: q <= 32'b10111101000010010101001011110010 ;
        2760: q <= 32'b00111101101110111000100100101100 ;
        2761: q <= 32'b10111100011000001100110001010100 ;
        2762: q <= 32'b10111101100001011100011111000011 ;
        2763: q <= 32'b00111101000010000111010011010111 ;
        2764: q <= 32'b00111100100011100110010000110111 ;
        2765: q <= 32'b00111100100110110100000100010111 ;
        2766: q <= 32'b00111100100110111011011011000011 ;
        2767: q <= 32'b00111100010110010101011000000100 ;
        2768: q <= 32'b00111011111000010100000001011100 ;
        2769: q <= 32'b00111101011101110001000100011000 ;
        2770: q <= 32'b10111110000000010001100100100010 ;
        2771: q <= 32'b10111110000011101010101010011000 ;
        2772: q <= 32'b10111100001011111111010000101000 ;
        2773: q <= 32'b10111011100110000001101010011011 ;
        2774: q <= 32'b00111101100011001100011011110100 ;
        2775: q <= 32'b10111101100101010101000101011110 ;
        2776: q <= 32'b10111100001111011101001000100100 ;
        2777: q <= 32'b10111101001101101111111010100000 ;
        2778: q <= 32'b10111101010110101111100101110100 ;
        2779: q <= 32'b10111101111100111111011000010000 ;
        2780: q <= 32'b00111100001100110101100101100100 ;
        2781: q <= 32'b00111100100011101101011001111100 ;
        2782: q <= 32'b10111101000000000000101111111110 ;
        2783: q <= 32'b10111100101010110010001001000000 ;
        2784: q <= 32'b00111101000101100011100001010011 ;
        2785: q <= 32'b10111101010101000110010110000011 ;
        2786: q <= 32'b10111100000010100100001001101000 ;
        2787: q <= 32'b10111110000001001000101100111110 ;
        2788: q <= 32'b00111100101001010010011000100011 ;
        2789: q <= 32'b00111101011001111011011000011110 ;
        2790: q <= 32'b10111100100110101010110001110010 ;
        2791: q <= 32'b10111101011110001001110001011001 ;
        2792: q <= 32'b00000000000000000000000000000000 ;
        2793: q <= 32'b00000000000000000000000000000000 ;
        2794: q <= 32'b00000000000000000000000000000000 ;
        2795: q <= 32'b00000000000000000000000000000000 ;
        2796: q <= 32'b00000000000000000000000000000000 ;
        2797: q <= 32'b00000000000000000000000000000000 ;
        2798: q <= 32'b00000000000000000000000000000000 ;
        2799: q <= 32'b00000000000000000000000000000000 ;
        2800: q <= 32'b00000000000000000000000000000000 ;
        2801: q <= 32'b00000000000000000000000000000000 ;
        2802: q <= 32'b00000000000000000000000000000000 ;
        2803: q <= 32'b00000000000000000000000000000000 ;
        2804: q <= 32'b00000000000000000000000000000000 ;
        2805: q <= 32'b00000000000000000000000000000000 ;
        2806: q <= 32'b00000000000000000000000000000000 ;
        2807: q <= 32'b00000000000000000000000000000000 ;
        2808: q <= 32'b00000000000000000000000000000000 ;
        2809: q <= 32'b00000000000000000000000000000000 ;
        2810: q <= 32'b00000000000000000000000000000000 ;
        2811: q <= 32'b00000000000000000000000000000000 ;
        2812: q <= 32'b00000000000000000000000000000000 ;
        2813: q <= 32'b00000000000000000000000000000000 ;
        2814: q <= 32'b00000000000000000000000000000000 ;
        2815: q <= 32'b00000000000000000000000000000000 ;
        2816: q <= 32'b10111101100001101010011111111101 ;
        2817: q <= 32'b00111110000011010100101000010000 ;
        2818: q <= 32'b10111101110100101100001001101001 ;
        2819: q <= 32'b00111100111000000111110010011000 ;
        2820: q <= 32'b00111110001101001010101101011111 ;
        2821: q <= 32'b10111101010001010111001100111100 ;
        2822: q <= 32'b10111101000010100110011000000110 ;
        2823: q <= 32'b00111101010000111101000100000001 ;
        2824: q <= 32'b10111110000000100010111000001110 ;
        2825: q <= 32'b00111101100110010001101011001011 ;
        2826: q <= 32'b00111101101011110110011111100101 ;
        2827: q <= 32'b00111101010010101110101101111001 ;
        2828: q <= 32'b10111101001110011001000111110111 ;
        2829: q <= 32'b00111011110010101111100011111100 ;
        2830: q <= 32'b00111101100110011010111001100110 ;
        2831: q <= 32'b10111101100000000011101011011111 ;
        2832: q <= 32'b10111100111001000111011101111011 ;
        2833: q <= 32'b10111101100011000010011000011110 ;
        2834: q <= 32'b10111011111011111000110101100110 ;
        2835: q <= 32'b00111101011010110001111100110000 ;
        2836: q <= 32'b10111101001111010010111001101111 ;
        2837: q <= 32'b10111101100000001001011101011011 ;
        2838: q <= 32'b00111100110101110000110011011000 ;
        2839: q <= 32'b00111101111101001011101000011010 ;
        2840: q <= 32'b00111101001001101011011111111010 ;
        2841: q <= 32'b00111101000011011000011001010000 ;
        2842: q <= 32'b10111101100001100100001000001101 ;
        2843: q <= 32'b00111110000000000000100001101111 ;
        2844: q <= 32'b10111101111000101011110100010001 ;
        2845: q <= 32'b10111101100000011000111111001011 ;
        2846: q <= 32'b00111110000011000000100100100001 ;
        2847: q <= 32'b10111101100000111110010000011010 ;
        2848: q <= 32'b10111101101100111110101000101110 ;
        2849: q <= 32'b00111100100111001001000000100010 ;
        2850: q <= 32'b10111101101110110010111001101000 ;
        2851: q <= 32'b00111011100001100110111001101110 ;
        2852: q <= 32'b00111101000001001001001111100101 ;
        2853: q <= 32'b10111101001110001010001000011100 ;
        2854: q <= 32'b10111100010110010010000111001001 ;
        2855: q <= 32'b00111100110011000100000001001100 ;
        2856: q <= 32'b00111101100010010010011010000110 ;
        2857: q <= 32'b10111101101101001001110011101111 ;
        2858: q <= 32'b00111100100110110001000111100010 ;
        2859: q <= 32'b10111101100001110100000011001110 ;
        2860: q <= 32'b00111101011001100010011010000101 ;
        2861: q <= 32'b00111011101100100101100101101000 ;
        2862: q <= 32'b10111101100001111100101100110110 ;
        2863: q <= 32'b00111101010111100010011001100110 ;
        2864: q <= 32'b10111101110110101101000111001001 ;
        2865: q <= 32'b00111101101001101110010101011101 ;
        2866: q <= 32'b10111100100110110000011101100111 ;
        2867: q <= 32'b00111101101010011000111011001110 ;
        2868: q <= 32'b00111100101101100011111010110011 ;
        2869: q <= 32'b00111101100111011111111100101110 ;
        2870: q <= 32'b10111101110101110101000101010001 ;
        2871: q <= 32'b00111100001110010101111100001010 ;
        2872: q <= 32'b00111101001001001010101001101101 ;
        2873: q <= 32'b10111011011110000100100110000011 ;
        2874: q <= 32'b10111101101011001100110011001010 ;
        2875: q <= 32'b00111100100011110101111110100110 ;
        2876: q <= 32'b00111101100101000100111101101111 ;
        2877: q <= 32'b00111100011110000000110001101100 ;
        2878: q <= 32'b00111100110110101000110101011010 ;
        2879: q <= 32'b10111100101111100001001100001111 ;
        2880: q <= 32'b10111101101110010101001000101101 ;
        2881: q <= 32'b10111101101101000010001001011010 ;
        2882: q <= 32'b00111101110101101110111001001001 ;
        2883: q <= 32'b10111100000010001000101111000110 ;
        2884: q <= 32'b00111110000000001110010110000111 ;
        2885: q <= 32'b00111101010111111100000000010101 ;
        2886: q <= 32'b00111100111010101111001110011111 ;
        2887: q <= 32'b00111100000010011001111001000010 ;
        2888: q <= 32'b10111100001101000101010011000001 ;
        2889: q <= 32'b10111101110011110000010110000010 ;
        2890: q <= 32'b00111101000011100111011100001001 ;
        2891: q <= 32'b10111101010101111110000011111110 ;
        2892: q <= 32'b10111101011101000001011010010000 ;
        2893: q <= 32'b00111101001111101110000111000000 ;
        2894: q <= 32'b00111100111010011101101000000010 ;
        2895: q <= 32'b00111101011111110101111111001011 ;
        2896: q <= 32'b10111110000001111110110101101111 ;
        2897: q <= 32'b00111101111110111011111101001101 ;
        2898: q <= 32'b00111100011100010010101110110010 ;
        2899: q <= 32'b10111101010110100101000000011101 ;
        2900: q <= 32'b00111100111011000001110000101111 ;
        2901: q <= 32'b10111100000101101010010000100101 ;
        2902: q <= 32'b00111011111111111111100101100010 ;
        2903: q <= 32'b00111101001110110101111100001110 ;
        2904: q <= 32'b00111101011111100000000010101110 ;
        2905: q <= 32'b00111101100010001001100100011100 ;
        2906: q <= 32'b10111101110001000010000010100101 ;
        2907: q <= 32'b00111101100110100101010110110111 ;
        2908: q <= 32'b10111101010001001100111011101000 ;
        2909: q <= 32'b10111101110100110010011010001010 ;
        2910: q <= 32'b00111101011010100010001010011001 ;
        2911: q <= 32'b10111101100101000000110110110001 ;
        2912: q <= 32'b00111110000011011000011011000000 ;
        2913: q <= 32'b00111101010000001111110100111110 ;
        2914: q <= 32'b10111101110000100111001011000010 ;
        2915: q <= 32'b00111101100101110111011011100010 ;
        2916: q <= 32'b10111011001001011111011110110100 ;
        2917: q <= 32'b00111100111111100111010011001000 ;
        2918: q <= 32'b10111100100110010111100000111000 ;
        2919: q <= 32'b10111100110100010111000100111010 ;
        2920: q <= 32'b00000000000000000000000000000000 ;
        2921: q <= 32'b00000000000000000000000000000000 ;
        2922: q <= 32'b00000000000000000000000000000000 ;
        2923: q <= 32'b00000000000000000000000000000000 ;
        2924: q <= 32'b00000000000000000000000000000000 ;
        2925: q <= 32'b00000000000000000000000000000000 ;
        2926: q <= 32'b00000000000000000000000000000000 ;
        2927: q <= 32'b00000000000000000000000000000000 ;
        2928: q <= 32'b00000000000000000000000000000000 ;
        2929: q <= 32'b00000000000000000000000000000000 ;
        2930: q <= 32'b00000000000000000000000000000000 ;
        2931: q <= 32'b00000000000000000000000000000000 ;
        2932: q <= 32'b00000000000000000000000000000000 ;
        2933: q <= 32'b00000000000000000000000000000000 ;
        2934: q <= 32'b00000000000000000000000000000000 ;
        2935: q <= 32'b00000000000000000000000000000000 ;
        2936: q <= 32'b00000000000000000000000000000000 ;
        2937: q <= 32'b00000000000000000000000000000000 ;
        2938: q <= 32'b00000000000000000000000000000000 ;
        2939: q <= 32'b00000000000000000000000000000000 ;
        2940: q <= 32'b00000000000000000000000000000000 ;
        2941: q <= 32'b00000000000000000000000000000000 ;
        2942: q <= 32'b00000000000000000000000000000000 ;
        2943: q <= 32'b00000000000000000000000000000000 ;
        2944: q <= 32'b00111101001101110111110111111010 ;
        2945: q <= 32'b10111100111000010010000101100110 ;
        2946: q <= 32'b00111101100010001011100000111001 ;
        2947: q <= 32'b00111101100010101111101010000100 ;
        2948: q <= 32'b10111101100111001000110000101101 ;
        2949: q <= 32'b00111101100000101010101110001001 ;
        2950: q <= 32'b00111101000011010100000000000101 ;
        2951: q <= 32'b10111100101101011001011001110101 ;
        2952: q <= 32'b10111101000001100110000110000111 ;
        2953: q <= 32'b00111101110011101111001000101100 ;
        2954: q <= 32'b10111110000000100110100001101100 ;
        2955: q <= 32'b00111110000111001010101011000000 ;
        2956: q <= 32'b00111101100110110000110000110011 ;
        2957: q <= 32'b00111101011010110001000111100101 ;
        2958: q <= 32'b10111100101101011010011010110000 ;
        2959: q <= 32'b00111100101100101100110010011110 ;
        2960: q <= 32'b00111101010010100110010111111001 ;
        2961: q <= 32'b10111101010101010001110100000011 ;
        2962: q <= 32'b00111101110010100000010001101010 ;
        2963: q <= 32'b10111100100000010010011011110000 ;
        2964: q <= 32'b10111101001100101010000100111100 ;
        2965: q <= 32'b00111110000110110100001101010101 ;
        2966: q <= 32'b10111100111100101101110010111010 ;
        2967: q <= 32'b10111101100000010000001110001001 ;
        2968: q <= 32'b10111101100001111100010001101101 ;
        2969: q <= 32'b10111011111100101011011110001011 ;
        2970: q <= 32'b00111101011101001000111011111010 ;
        2971: q <= 32'b10111011110111000010000101010111 ;
        2972: q <= 32'b00111100101010001010111100011100 ;
        2973: q <= 32'b10111101000001101110100001000001 ;
        2974: q <= 32'b00111101101100111011111000001010 ;
        2975: q <= 32'b10111100110110111100011001110101 ;
        2976: q <= 32'b10111101101000111010110001110111 ;
        2977: q <= 32'b00111101101001001001010011101100 ;
        2978: q <= 32'b00111101100010100000001111010000 ;
        2979: q <= 32'b00111110000000000010010010000000 ;
        2980: q <= 32'b10111101111100010001000010000000 ;
        2981: q <= 32'b10111100000101110101001010000101 ;
        2982: q <= 32'b10111101100000010100001110100000 ;
        2983: q <= 32'b00111101000011100000101101000000 ;
        2984: q <= 32'b10111101101000010101000110101010 ;
        2985: q <= 32'b00111101001111000110011111111111 ;
        2986: q <= 32'b10111100010110010111100110101010 ;
        2987: q <= 32'b00111100001111111000100001110100 ;
        2988: q <= 32'b00111100101010111010010000011111 ;
        2989: q <= 32'b00111101100001000111100110001011 ;
        2990: q <= 32'b10111101010101011001100011110000 ;
        2991: q <= 32'b00111101111011001101101111111110 ;
        2992: q <= 32'b00111101001000011111000100101001 ;
        2993: q <= 32'b00111101100100010011101110100000 ;
        2994: q <= 32'b10111101100100111001010011111111 ;
        2995: q <= 32'b10111100000101010110100101011001 ;
        2996: q <= 32'b10111101101000101101000100010001 ;
        2997: q <= 32'b10111101101010011010100110111011 ;
        2998: q <= 32'b00111101101101110001100111101000 ;
        2999: q <= 32'b10111101011000100010011011100100 ;
        3000: q <= 32'b00111101110010101101000100001001 ;
        3001: q <= 32'b10111101111011101000001100000100 ;
        3002: q <= 32'b10111101101100110100110000111000 ;
        3003: q <= 32'b00111101101001111010110100010001 ;
        3004: q <= 32'b10111100001100111000101100000111 ;
        3005: q <= 32'b10111100111001100100110001100011 ;
        3006: q <= 32'b00111100110001110010001110110000 ;
        3007: q <= 32'b00111101010101011100010010000111 ;
        3008: q <= 32'b00111010011010011111000000001010 ;
        3009: q <= 32'b10111100000110111111111101010011 ;
        3010: q <= 32'b00111100101000111110001111010110 ;
        3011: q <= 32'b00111101011011101011111101011111 ;
        3012: q <= 32'b10111101001011111110001011111000 ;
        3013: q <= 32'b10111100111010100000011011001111 ;
        3014: q <= 32'b10111100100011110000101100111101 ;
        3015: q <= 32'b10111110000100001100010110001000 ;
        3016: q <= 32'b10111100110100000111100100010100 ;
        3017: q <= 32'b10111010000111101110011111010000 ;
        3018: q <= 32'b00111101001010010101101010011011 ;
        3019: q <= 32'b00111110000100101011010000100100 ;
        3020: q <= 32'b10111110000010101101011101001111 ;
        3021: q <= 32'b00111101100011100100111011100001 ;
        3022: q <= 32'b10111101011010101010110010111010 ;
        3023: q <= 32'b00111101110101011010010011000001 ;
        3024: q <= 32'b00111101111001110011010110101101 ;
        3025: q <= 32'b10111101101110101000001101011010 ;
        3026: q <= 32'b00111101000011000010001000001111 ;
        3027: q <= 32'b00111101101100101001010011000001 ;
        3028: q <= 32'b10111110000111101111001000111110 ;
        3029: q <= 32'b00111100111101001001100101101111 ;
        3030: q <= 32'b10111101000101000110001001010101 ;
        3031: q <= 32'b00111101101110110110011111011000 ;
        3032: q <= 32'b10111101011100101011011010110110 ;
        3033: q <= 32'b10111101100001111011110111001110 ;
        3034: q <= 32'b10111101100010111011110010110011 ;
        3035: q <= 32'b10111100110101010001101100011110 ;
        3036: q <= 32'b00111101100100010100000100100001 ;
        3037: q <= 32'b00111101111001101110101111000101 ;
        3038: q <= 32'b00111101110100000101010100111101 ;
        3039: q <= 32'b00111101011000111100100110010010 ;
        3040: q <= 32'b00111101010111010011001000101101 ;
        3041: q <= 32'b00111100001010001110010110110111 ;
        3042: q <= 32'b10111100111001111010111000100011 ;
        3043: q <= 32'b00111101100111011110111110101010 ;
        3044: q <= 32'b00111101100011000000011000010010 ;
        3045: q <= 32'b00111100101010101101011010100001 ;
        3046: q <= 32'b10111101100100100101000010111100 ;
        3047: q <= 32'b10111101100000111000101101111011 ;
        3048: q <= 32'b00000000000000000000000000000000 ;
        3049: q <= 32'b00000000000000000000000000000000 ;
        3050: q <= 32'b00000000000000000000000000000000 ;
        3051: q <= 32'b00000000000000000000000000000000 ;
        3052: q <= 32'b00000000000000000000000000000000 ;
        3053: q <= 32'b00000000000000000000000000000000 ;
        3054: q <= 32'b00000000000000000000000000000000 ;
        3055: q <= 32'b00000000000000000000000000000000 ;
        3056: q <= 32'b00000000000000000000000000000000 ;
        3057: q <= 32'b00000000000000000000000000000000 ;
        3058: q <= 32'b00000000000000000000000000000000 ;
        3059: q <= 32'b00000000000000000000000000000000 ;
        3060: q <= 32'b00000000000000000000000000000000 ;
        3061: q <= 32'b00000000000000000000000000000000 ;
        3062: q <= 32'b00000000000000000000000000000000 ;
        3063: q <= 32'b00000000000000000000000000000000 ;
        3064: q <= 32'b00000000000000000000000000000000 ;
        3065: q <= 32'b00000000000000000000000000000000 ;
        3066: q <= 32'b00000000000000000000000000000000 ;
        3067: q <= 32'b00000000000000000000000000000000 ;
        3068: q <= 32'b00000000000000000000000000000000 ;
        3069: q <= 32'b00000000000000000000000000000000 ;
        3070: q <= 32'b00000000000000000000000000000000 ;
        3071: q <= 32'b00000000000000000000000000000000 ;
        3072: q <= 32'b00111101110010011010010111010110 ;
        3073: q <= 32'b00111100111110001011010110101011 ;
        3074: q <= 32'b00111011101110101101110100011001 ;
        3075: q <= 32'b00111101000111110101110110101010 ;
        3076: q <= 32'b00111100110110110110011111111111 ;
        3077: q <= 32'b00111101100000001010100001010111 ;
        3078: q <= 32'b00111101000110001101100100001001 ;
        3079: q <= 32'b10111101100000111011100000000100 ;
        3080: q <= 32'b10111101101000100111110111001010 ;
        3081: q <= 32'b00111101011000110000000010010000 ;
        3082: q <= 32'b00111100111101101110100111111011 ;
        3083: q <= 32'b00111101101100000111111111111110 ;
        3084: q <= 32'b10111100011001101110010111001111 ;
        3085: q <= 32'b00111101001001000000101110101000 ;
        3086: q <= 32'b00111100001101010010110110001001 ;
        3087: q <= 32'b00111101011110000110001000110101 ;
        3088: q <= 32'b00111101011011000001001100101110 ;
        3089: q <= 32'b00111101110101001110010110010001 ;
        3090: q <= 32'b00111110001100011011111100001110 ;
        3091: q <= 32'b10111110000110111011101101101011 ;
        3092: q <= 32'b10111101001110100000010001000000 ;
        3093: q <= 32'b00111101101001010001111001001010 ;
        3094: q <= 32'b10111101111000001000110000001101 ;
        3095: q <= 32'b10111101011001001011110100000110 ;
        3096: q <= 32'b10111101001110000000000010101110 ;
        3097: q <= 32'b10111110000010010001011010000111 ;
        3098: q <= 32'b00111100111010011010001011110111 ;
        3099: q <= 32'b00111011001011110100110100110010 ;
        3100: q <= 32'b00111100100111101001011100110110 ;
        3101: q <= 32'b00111101101111000000111000100111 ;
        3102: q <= 32'b00111110001010101010101000111110 ;
        3103: q <= 32'b10111101001010101011111000011111 ;
        3104: q <= 32'b00111100100011011001111100111011 ;
        3105: q <= 32'b00111011011110111001001011111010 ;
        3106: q <= 32'b00111101001101001011110100010110 ;
        3107: q <= 32'b10111101010011101011101101001110 ;
        3108: q <= 32'b10111101101110111010101000101001 ;
        3109: q <= 32'b00111110000010011001100111110011 ;
        3110: q <= 32'b00111100001000011101010000100110 ;
        3111: q <= 32'b00111101110100010100001111111011 ;
        3112: q <= 32'b10111101010100111001111100100011 ;
        3113: q <= 32'b00111101100101101000111100111000 ;
        3114: q <= 32'b00111101011100111101100101011000 ;
        3115: q <= 32'b10111110000011011010000110110101 ;
        3116: q <= 32'b10111101100001000101000110110001 ;
        3117: q <= 32'b10111101101111111000110011110101 ;
        3118: q <= 32'b00111101110001100011010110101011 ;
        3119: q <= 32'b00111101001011001101000001110101 ;
        3120: q <= 32'b00111011000111100001010001101101 ;
        3121: q <= 32'b00111101000011110001011100001101 ;
        3122: q <= 32'b00111100110000111000110001111010 ;
        3123: q <= 32'b10111101010011100001111011010001 ;
        3124: q <= 32'b10111101100100110001101000010111 ;
        3125: q <= 32'b10111110000000101111010000011101 ;
        3126: q <= 32'b00111110010010010000001000111101 ;
        3127: q <= 32'b00111101010100110001011101011011 ;
        3128: q <= 32'b00111101111110010011110001110101 ;
        3129: q <= 32'b10111101010100011101111110001111 ;
        3130: q <= 32'b10111101110011111111111001000010 ;
        3131: q <= 32'b10111101011110000011001010011111 ;
        3132: q <= 32'b10111100011011100001100110101011 ;
        3133: q <= 32'b00111100111010110110010000000111 ;
        3134: q <= 32'b10111101000010000011101100111001 ;
        3135: q <= 32'b00111101101110000011111011001001 ;
        3136: q <= 32'b00111101101110110101111011111001 ;
        3137: q <= 32'b00111011100010111010100000101101 ;
        3138: q <= 32'b10111101100000101100100101010100 ;
        3139: q <= 32'b00111101000000110111101101010001 ;
        3140: q <= 32'b10111101100110011101010111010100 ;
        3141: q <= 32'b10111100000000000000010111111000 ;
        3142: q <= 32'b10111011010000110000000011011010 ;
        3143: q <= 32'b10111110000110011010011100111101 ;
        3144: q <= 32'b10111100100101101101100100110000 ;
        3145: q <= 32'b10111101100011011011010110100110 ;
        3146: q <= 32'b00111101001011000100001010110110 ;
        3147: q <= 32'b00111101001011100001110011111011 ;
        3148: q <= 32'b10111110000101001111001001110100 ;
        3149: q <= 32'b10111000111000000001000110110010 ;
        3150: q <= 32'b10111101100111001010000111010000 ;
        3151: q <= 32'b00111110000000111010110000011100 ;
        3152: q <= 32'b10111101110000011010100100011101 ;
        3153: q <= 32'b10111101110100111111011111101001 ;
        3154: q <= 32'b00111110001000001001101010000000 ;
        3155: q <= 32'b00111101100110010011110111100111 ;
        3156: q <= 32'b10111110000000010100100100011001 ;
        3157: q <= 32'b10111100101110011011011111111110 ;
        3158: q <= 32'b00111100111001111100011001001111 ;
        3159: q <= 32'b10111101100000111111101111100010 ;
        3160: q <= 32'b10111101101100101110100111000001 ;
        3161: q <= 32'b00111100110001101000111100000000 ;
        3162: q <= 32'b10111100100010001101010000000001 ;
        3163: q <= 32'b10111100110010100100011000111000 ;
        3164: q <= 32'b10111101101011010100110101000001 ;
        3165: q <= 32'b00111101100011111101001000111100 ;
        3166: q <= 32'b10111101011101001010010000101111 ;
        3167: q <= 32'b00111101110000101101101101110111 ;
        3168: q <= 32'b00111101011001111111111000011010 ;
        3169: q <= 32'b00111100100111011100101001100111 ;
        3170: q <= 32'b00111101110110000001100001111111 ;
        3171: q <= 32'b10111101001111110000101101001011 ;
        3172: q <= 32'b10111101010011000010111100101001 ;
        3173: q <= 32'b00111101011100101110011101100000 ;
        3174: q <= 32'b00111101000000110101110011000100 ;
        3175: q <= 32'b00111101101011110000101100111101 ;
        3176: q <= 32'b00000000000000000000000000000000 ;
        3177: q <= 32'b00000000000000000000000000000000 ;
        3178: q <= 32'b00000000000000000000000000000000 ;
        3179: q <= 32'b00000000000000000000000000000000 ;
        3180: q <= 32'b00000000000000000000000000000000 ;
        3181: q <= 32'b00000000000000000000000000000000 ;
        3182: q <= 32'b00000000000000000000000000000000 ;
        3183: q <= 32'b00000000000000000000000000000000 ;
        3184: q <= 32'b00000000000000000000000000000000 ;
        3185: q <= 32'b00000000000000000000000000000000 ;
        3186: q <= 32'b00000000000000000000000000000000 ;
        3187: q <= 32'b00000000000000000000000000000000 ;
        3188: q <= 32'b00000000000000000000000000000000 ;
        3189: q <= 32'b00000000000000000000000000000000 ;
        3190: q <= 32'b00000000000000000000000000000000 ;
        3191: q <= 32'b00000000000000000000000000000000 ;
        3192: q <= 32'b00000000000000000000000000000000 ;
        3193: q <= 32'b00000000000000000000000000000000 ;
        3194: q <= 32'b00000000000000000000000000000000 ;
        3195: q <= 32'b00000000000000000000000000000000 ;
        3196: q <= 32'b00000000000000000000000000000000 ;
        3197: q <= 32'b00000000000000000000000000000000 ;
        3198: q <= 32'b00000000000000000000000000000000 ;
        3199: q <= 32'b00000000000000000000000000000000 ;
        3200: q <= 32'b10111101110101111100101100110110 ;
        3201: q <= 32'b00111101100000010100101000001110 ;
        3202: q <= 32'b10111110000011001100110010110001 ;
        3203: q <= 32'b00111100000000000010010101101011 ;
        3204: q <= 32'b00111101011101111101000100111110 ;
        3205: q <= 32'b00111101000110110101001011011100 ;
        3206: q <= 32'b10111101100010101000011110101100 ;
        3207: q <= 32'b00111100010010110111101000101110 ;
        3208: q <= 32'b00111101100001010110000010010010 ;
        3209: q <= 32'b10111010001010001111000010011001 ;
        3210: q <= 32'b10111100111101000001011010001111 ;
        3211: q <= 32'b10111101101111011001100000101010 ;
        3212: q <= 32'b00111101101011001110100001101110 ;
        3213: q <= 32'b00111100011000010110011000010101 ;
        3214: q <= 32'b10111101000100001110110100100110 ;
        3215: q <= 32'b10111011111110001010000100100000 ;
        3216: q <= 32'b10111011100011110011000011011111 ;
        3217: q <= 32'b10111101101001111100101110110001 ;
        3218: q <= 32'b10111101100101111101100100100111 ;
        3219: q <= 32'b10111101001001100111100000000101 ;
        3220: q <= 32'b00111101101111001101010111001000 ;
        3221: q <= 32'b10111101100100010001000111001100 ;
        3222: q <= 32'b10111101010000001110010111001000 ;
        3223: q <= 32'b00111100010010000001100111010001 ;
        3224: q <= 32'b00111100011000100011011111101010 ;
        3225: q <= 32'b10111101100011100011011001110101 ;
        3226: q <= 32'b10111101000000001000001000111000 ;
        3227: q <= 32'b10111101101100110100000010010101 ;
        3228: q <= 32'b10111101000100101001111101111111 ;
        3229: q <= 32'b00111101011100010001110001001001 ;
        3230: q <= 32'b10111011001100010010111001010001 ;
        3231: q <= 32'b10111101101000000001010000000111 ;
        3232: q <= 32'b00111011100011111001010100001011 ;
        3233: q <= 32'b00111101101100111010010111011011 ;
        3234: q <= 32'b10111101011101001101001011011100 ;
        3235: q <= 32'b10111100111001111010010100001101 ;
        3236: q <= 32'b10111101010000000111011101101010 ;
        3237: q <= 32'b00111101101100010010111001110010 ;
        3238: q <= 32'b00111101011110010001110001010101 ;
        3239: q <= 32'b00111011110000111000011111110110 ;
        3240: q <= 32'b10111101011101010001010010111010 ;
        3241: q <= 32'b10111101011100001110101011001001 ;
        3242: q <= 32'b00111100011011011001010001110101 ;
        3243: q <= 32'b10111101100010010001111010110101 ;
        3244: q <= 32'b10111101010110100001110101000010 ;
        3245: q <= 32'b10111100001100111010001011100010 ;
        3246: q <= 32'b00111101101011010010111001101100 ;
        3247: q <= 32'b10111101101010011010010100011001 ;
        3248: q <= 32'b10111100001111111101000011000011 ;
        3249: q <= 32'b00111101100010100110111100100100 ;
        3250: q <= 32'b00111101101010000011101111010011 ;
        3251: q <= 32'b00111101000001110011011001101011 ;
        3252: q <= 32'b10111101111100010111110001111110 ;
        3253: q <= 32'b00111101001000011110000011101011 ;
        3254: q <= 32'b10111100001100011100101101001001 ;
        3255: q <= 32'b10111100001101011100011001011111 ;
        3256: q <= 32'b10111101101001010110000010100011 ;
        3257: q <= 32'b00111101100111110001001001110000 ;
        3258: q <= 32'b10111101010100100110100000011100 ;
        3259: q <= 32'b00111101001110010111110111011001 ;
        3260: q <= 32'b00111101110001000101111110010010 ;
        3261: q <= 32'b10111101010001010101100100001011 ;
        3262: q <= 32'b10111100110110010010010001100101 ;
        3263: q <= 32'b10111101101101110110100101111000 ;
        3264: q <= 32'b10111101011101101100100100011011 ;
        3265: q <= 32'b00111011101111001111110111100101 ;
        3266: q <= 32'b00111100001101100011001010110111 ;
        3267: q <= 32'b10111100000000001111110100110110 ;
        3268: q <= 32'b00111100111110000000011000100110 ;
        3269: q <= 32'b00111101100100110000110010011100 ;
        3270: q <= 32'b00111101001011000101011001100101 ;
        3271: q <= 32'b00111100110100010010011011010010 ;
        3272: q <= 32'b10111101001001000100001010011100 ;
        3273: q <= 32'b00111101011110001001011011100101 ;
        3274: q <= 32'b00111100010000110011011000111110 ;
        3275: q <= 32'b00111101011011000100100011011000 ;
        3276: q <= 32'b00111100101101000101110111010110 ;
        3277: q <= 32'b00111100000111101011101011100100 ;
        3278: q <= 32'b10111100101100011011101101010000 ;
        3279: q <= 32'b10111101100110000010111111001100 ;
        3280: q <= 32'b10111101100100011000011001001110 ;
        3281: q <= 32'b00111100101011001110000111111101 ;
        3282: q <= 32'b10111101011010001100111001110101 ;
        3283: q <= 32'b10111011101110011111010000010011 ;
        3284: q <= 32'b10111101000101111001110100011110 ;
        3285: q <= 32'b00111101010110100111110001011011 ;
        3286: q <= 32'b10111101101000110001111010001100 ;
        3287: q <= 32'b00111101000010001111001111100110 ;
        3288: q <= 32'b10111101100000101000110001011101 ;
        3289: q <= 32'b00111100111101111110110110101000 ;
        3290: q <= 32'b10111100110110110110101100011000 ;
        3291: q <= 32'b10111011101110011010000100001111 ;
        3292: q <= 32'b00111101100110101010001110000001 ;
        3293: q <= 32'b10111011111001111101000001011110 ;
        3294: q <= 32'b10111101101011101101010011111011 ;
        3295: q <= 32'b10111011110001010011011111101111 ;
        3296: q <= 32'b10111101100000111100010011000001 ;
        3297: q <= 32'b00111100100100001000110110101011 ;
        3298: q <= 32'b00111101010100011000011011100100 ;
        3299: q <= 32'b00111101010001001100111001010011 ;
        3300: q <= 32'b00111011001100101010011110000010 ;
        3301: q <= 32'b10111101000101101000110001000111 ;
        3302: q <= 32'b10111100000011111100000001011100 ;
        3303: q <= 32'b10111101110001010100011101000011 ;
        3304: q <= 32'b00000000000000000000000000000000 ;
        3305: q <= 32'b00000000000000000000000000000000 ;
        3306: q <= 32'b00000000000000000000000000000000 ;
        3307: q <= 32'b00000000000000000000000000000000 ;
        3308: q <= 32'b00000000000000000000000000000000 ;
        3309: q <= 32'b00000000000000000000000000000000 ;
        3310: q <= 32'b00000000000000000000000000000000 ;
        3311: q <= 32'b00000000000000000000000000000000 ;
        3312: q <= 32'b00000000000000000000000000000000 ;
        3313: q <= 32'b00000000000000000000000000000000 ;
        3314: q <= 32'b00000000000000000000000000000000 ;
        3315: q <= 32'b00000000000000000000000000000000 ;
        3316: q <= 32'b00000000000000000000000000000000 ;
        3317: q <= 32'b00000000000000000000000000000000 ;
        3318: q <= 32'b00000000000000000000000000000000 ;
        3319: q <= 32'b00000000000000000000000000000000 ;
        3320: q <= 32'b00000000000000000000000000000000 ;
        3321: q <= 32'b00000000000000000000000000000000 ;
        3322: q <= 32'b00000000000000000000000000000000 ;
        3323: q <= 32'b00000000000000000000000000000000 ;
        3324: q <= 32'b00000000000000000000000000000000 ;
        3325: q <= 32'b00000000000000000000000000000000 ;
        3326: q <= 32'b00000000000000000000000000000000 ;
        3327: q <= 32'b00000000000000000000000000000000 ;
        3328: q <= 32'b00111011111000011000010011101010 ;
        3329: q <= 32'b00111011100001010010001000101010 ;
        3330: q <= 32'b00111100100011110011111001000101 ;
        3331: q <= 32'b10111101011010111110000111101010 ;
        3332: q <= 32'b10111101001110110011111010001000 ;
        3333: q <= 32'b00111101000101101110010100000001 ;
        3334: q <= 32'b10111101110000110000110101100011 ;
        3335: q <= 32'b10111101010011000100011100100110 ;
        3336: q <= 32'b00111101111001111101110011111001 ;
        3337: q <= 32'b10111010010111111011010100011111 ;
        3338: q <= 32'b10111101100011011000011101101101 ;
        3339: q <= 32'b00111100101111110000010110110100 ;
        3340: q <= 32'b10111101110100011001111000010001 ;
        3341: q <= 32'b00111110001001111001001011111010 ;
        3342: q <= 32'b10111101110110101111101001101100 ;
        3343: q <= 32'b00111100101111110001010001010001 ;
        3344: q <= 32'b00111110000000000001110001101001 ;
        3345: q <= 32'b00111101111100101110010111001110 ;
        3346: q <= 32'b10111011100111000100011111010110 ;
        3347: q <= 32'b10111110011111101100100101111110 ;
        3348: q <= 32'b00111100000010111110011110111100 ;
        3349: q <= 32'b10111101101011001001001111111111 ;
        3350: q <= 32'b00111110010110101010110100011110 ;
        3351: q <= 32'b00111100111011011110101000111000 ;
        3352: q <= 32'b10111101101101110111100010011010 ;
        3353: q <= 32'b10111101010100000100100001110110 ;
        3354: q <= 32'b10111100001010111011111101101100 ;
        3355: q <= 32'b10111101000000111111110010011111 ;
        3356: q <= 32'b10111100101011101110110110000100 ;
        3357: q <= 32'b00111101010010101001001111101001 ;
        3358: q <= 32'b10111011101100000010100101100100 ;
        3359: q <= 32'b00111100101011100101001110011011 ;
        3360: q <= 32'b00111100101110101101101111101110 ;
        3361: q <= 32'b10111101011101100000100010000001 ;
        3362: q <= 32'b10111101010010110111011110101001 ;
        3363: q <= 32'b10111011110111110101011111001110 ;
        3364: q <= 32'b00111101100001000010001110101110 ;
        3365: q <= 32'b00111101100001110011000000001010 ;
        3366: q <= 32'b10111101101010000111100010110110 ;
        3367: q <= 32'b00111101111100100001011101110011 ;
        3368: q <= 32'b10111011010110101001001010111101 ;
        3369: q <= 32'b10111101100010001001101000101111 ;
        3370: q <= 32'b00111101100011000101011011100000 ;
        3371: q <= 32'b00111101000110000000111111011111 ;
        3372: q <= 32'b10111110001100111100001101000100 ;
        3373: q <= 32'b00111101001110111110100110101000 ;
        3374: q <= 32'b10111101011001101001101001011100 ;
        3375: q <= 32'b10111101100011001110010111110000 ;
        3376: q <= 32'b00111101101011011010100010100010 ;
        3377: q <= 32'b10111101011100110100101000011101 ;
        3378: q <= 32'b00111101100110111100011111100101 ;
        3379: q <= 32'b00111100100101101011100000110100 ;
        3380: q <= 32'b00111101111110110000101001000010 ;
        3381: q <= 32'b00111101111011110101010100111101 ;
        3382: q <= 32'b10111100101001010100001110011110 ;
        3383: q <= 32'b00111101101101100110001110000101 ;
        3384: q <= 32'b00111101001111010101110101110101 ;
        3385: q <= 32'b10111011001101111110111101111111 ;
        3386: q <= 32'b10111101110000011100000101001110 ;
        3387: q <= 32'b10111101100011000001100111010111 ;
        3388: q <= 32'b10111101110000001101100101101001 ;
        3389: q <= 32'b10111100100111100100101111011000 ;
        3390: q <= 32'b00111101000010000111101011110110 ;
        3391: q <= 32'b00111101101010001101000101110010 ;
        3392: q <= 32'b10111101100100010110101011101001 ;
        3393: q <= 32'b00111101011010101001111111010000 ;
        3394: q <= 32'b00111101011111100101001001111101 ;
        3395: q <= 32'b10111101101110100110101111011100 ;
        3396: q <= 32'b00111101011011110101001101110000 ;
        3397: q <= 32'b10111101100001001101110010111000 ;
        3398: q <= 32'b10111101110110011011101100100101 ;
        3399: q <= 32'b10111100111011111110110011001100 ;
        3400: q <= 32'b10111100001100101000000000010100 ;
        3401: q <= 32'b10111011101111011011011000110110 ;
        3402: q <= 32'b10111011111010001011111111110110 ;
        3403: q <= 32'b00111101001000000011100010110100 ;
        3404: q <= 32'b00111101100001011001110101101111 ;
        3405: q <= 32'b10111101101011010111011110100010 ;
        3406: q <= 32'b10111101010101011101000100010001 ;
        3407: q <= 32'b00111100111101000011111000011100 ;
        3408: q <= 32'b10111101010001010101001100010111 ;
        3409: q <= 32'b00111101001101101101010001101011 ;
        3410: q <= 32'b00111110000000001100001011100011 ;
        3411: q <= 32'b10111100111011011010110011011100 ;
        3412: q <= 32'b10111101001100000110001101101010 ;
        3413: q <= 32'b00111100000010011011111011100000 ;
        3414: q <= 32'b00111101010010000000110101110000 ;
        3415: q <= 32'b00111101001110010111110110111110 ;
        3416: q <= 32'b00111101001101101100000011000100 ;
        3417: q <= 32'b10111101100101110101111110010100 ;
        3418: q <= 32'b00111101100100010100011110000111 ;
        3419: q <= 32'b00111101001110001110010111110010 ;
        3420: q <= 32'b10111100010101001110010011011101 ;
        3421: q <= 32'b10111100010011010111100110001111 ;
        3422: q <= 32'b10111100101111111000101001110111 ;
        3423: q <= 32'b00111101010100000110001000000110 ;
        3424: q <= 32'b10111101100100001100000101101111 ;
        3425: q <= 32'b00111101100110111101100100011001 ;
        3426: q <= 32'b00111110001000100011101001111110 ;
        3427: q <= 32'b00111101001110001110000001111000 ;
        3428: q <= 32'b10111011010011101101011001010000 ;
        3429: q <= 32'b00111100000111001001111111010110 ;
        3430: q <= 32'b00111101000001000110110101101000 ;
        3431: q <= 32'b10111101011101010110110101111101 ;
        3432: q <= 32'b00000000000000000000000000000000 ;
        3433: q <= 32'b00000000000000000000000000000000 ;
        3434: q <= 32'b00000000000000000000000000000000 ;
        3435: q <= 32'b00000000000000000000000000000000 ;
        3436: q <= 32'b00000000000000000000000000000000 ;
        3437: q <= 32'b00000000000000000000000000000000 ;
        3438: q <= 32'b00000000000000000000000000000000 ;
        3439: q <= 32'b00000000000000000000000000000000 ;
        3440: q <= 32'b00000000000000000000000000000000 ;
        3441: q <= 32'b00000000000000000000000000000000 ;
        3442: q <= 32'b00000000000000000000000000000000 ;
        3443: q <= 32'b00000000000000000000000000000000 ;
        3444: q <= 32'b00000000000000000000000000000000 ;
        3445: q <= 32'b00000000000000000000000000000000 ;
        3446: q <= 32'b00000000000000000000000000000000 ;
        3447: q <= 32'b00000000000000000000000000000000 ;
        3448: q <= 32'b00000000000000000000000000000000 ;
        3449: q <= 32'b00000000000000000000000000000000 ;
        3450: q <= 32'b00000000000000000000000000000000 ;
        3451: q <= 32'b00000000000000000000000000000000 ;
        3452: q <= 32'b00000000000000000000000000000000 ;
        3453: q <= 32'b00000000000000000000000000000000 ;
        3454: q <= 32'b00000000000000000000000000000000 ;
        3455: q <= 32'b00000000000000000000000000000000 ;
        3456: q <= 32'b00111100001010000010000101110000 ;
        3457: q <= 32'b10111100101001101101000111111010 ;
        3458: q <= 32'b10111101010010000111100100010001 ;
        3459: q <= 32'b10111101110000001010001001111010 ;
        3460: q <= 32'b10111101110001011111100100000101 ;
        3461: q <= 32'b10111101110100010101011000111100 ;
        3462: q <= 32'b10111101001000111001010000000110 ;
        3463: q <= 32'b10111101110010111011101010111000 ;
        3464: q <= 32'b00111101010110100011000011000100 ;
        3465: q <= 32'b00111101011101011001011110100010 ;
        3466: q <= 32'b10111101011101011001010100010100 ;
        3467: q <= 32'b00111101100110100000011100001100 ;
        3468: q <= 32'b00111101100010100000101101110101 ;
        3469: q <= 32'b00111100101000000000010111110001 ;
        3470: q <= 32'b00111100100011011110000101110010 ;
        3471: q <= 32'b10111011001110000111001011100110 ;
        3472: q <= 32'b10111100011101111110100110000111 ;
        3473: q <= 32'b00111101000101001011000100110000 ;
        3474: q <= 32'b10111011000111001100111000001110 ;
        3475: q <= 32'b10111101110000111110010000111011 ;
        3476: q <= 32'b10111100111110000000000000001111 ;
        3477: q <= 32'b00111101101110111011000110000110 ;
        3478: q <= 32'b10111011001101011011110011111001 ;
        3479: q <= 32'b10111101000101111110110000111101 ;
        3480: q <= 32'b00111100110111011111010100010101 ;
        3481: q <= 32'b10111100111100011010010010101100 ;
        3482: q <= 32'b10111110000010000101110011011100 ;
        3483: q <= 32'b10111101010101011011111011101001 ;
        3484: q <= 32'b10111101000001111011101111110110 ;
        3485: q <= 32'b10111010101101100000111010111000 ;
        3486: q <= 32'b10111101100000000101000100100110 ;
        3487: q <= 32'b00111101100011011000101111011001 ;
        3488: q <= 32'b00111101010101010100011010100111 ;
        3489: q <= 32'b10111101110000011110110000100001 ;
        3490: q <= 32'b00111101100011100110100100010000 ;
        3491: q <= 32'b10111101100111110101101110110100 ;
        3492: q <= 32'b00111101000001101000010010111101 ;
        3493: q <= 32'b10111101010111010110100100111010 ;
        3494: q <= 32'b00111101100101000011011100111110 ;
        3495: q <= 32'b00111101001010100111011111010011 ;
        3496: q <= 32'b10111101011100100001110100000011 ;
        3497: q <= 32'b10111100110001100011100100001000 ;
        3498: q <= 32'b00111101101111100000101110000101 ;
        3499: q <= 32'b00111011111100110000001110000011 ;
        3500: q <= 32'b00111101001000010110010100101101 ;
        3501: q <= 32'b00111101110001111100111101011110 ;
        3502: q <= 32'b10111101010001101100011000100011 ;
        3503: q <= 32'b00111101011110100101110000110100 ;
        3504: q <= 32'b10111001011010010111111000000110 ;
        3505: q <= 32'b00111101101000000011001101111100 ;
        3506: q <= 32'b10111101100101100101000001001111 ;
        3507: q <= 32'b00111100101101100000011110000111 ;
        3508: q <= 32'b10111100101011011110101001110111 ;
        3509: q <= 32'b00111100101101010111000001011101 ;
        3510: q <= 32'b10111100101011000010010011101011 ;
        3511: q <= 32'b10111101000000111000001101101011 ;
        3512: q <= 32'b00111101001000000010110000101011 ;
        3513: q <= 32'b00111101001101100011010010101101 ;
        3514: q <= 32'b00111101100110100011110001110000 ;
        3515: q <= 32'b10111101001110001101111111001110 ;
        3516: q <= 32'b00111101000010001101011001001011 ;
        3517: q <= 32'b10111101110001011000010010110011 ;
        3518: q <= 32'b10111101000000010001001001101111 ;
        3519: q <= 32'b00111100000001100000011011001101 ;
        3520: q <= 32'b00111101100111001111010011010100 ;
        3521: q <= 32'b00111101101110110111010010100010 ;
        3522: q <= 32'b00111101011011110100100010000010 ;
        3523: q <= 32'b00111101001101100110011101101001 ;
        3524: q <= 32'b10111100011001111100001001110111 ;
        3525: q <= 32'b00111100110011101111011010100001 ;
        3526: q <= 32'b00111101101000101101110000011001 ;
        3527: q <= 32'b00111101011111011110101100101110 ;
        3528: q <= 32'b10111101101010101001101101011001 ;
        3529: q <= 32'b10111101100111110111110010000001 ;
        3530: q <= 32'b10111101100100000011010011001111 ;
        3531: q <= 32'b00111011010000101010100001010001 ;
        3532: q <= 32'b00111101100110111000110001000111 ;
        3533: q <= 32'b10111100100011100111111001001101 ;
        3534: q <= 32'b10111101110011101001000110001100 ;
        3535: q <= 32'b10111101000111110110011111011000 ;
        3536: q <= 32'b10111101000000100101101111101100 ;
        3537: q <= 32'b00111101100100011101111001101011 ;
        3538: q <= 32'b00111101010100100011000001000111 ;
        3539: q <= 32'b00111101011010101110010011100001 ;
        3540: q <= 32'b00111101000100101101011101000110 ;
        3541: q <= 32'b00111101100001010011010010100111 ;
        3542: q <= 32'b10111101010000000011101001101001 ;
        3543: q <= 32'b10111101010000001001000111000001 ;
        3544: q <= 32'b10111101110010101010100111101000 ;
        3545: q <= 32'b00111101001011000011011111111001 ;
        3546: q <= 32'b00111100011010000000000100010011 ;
        3547: q <= 32'b10111101011001010111001100110100 ;
        3548: q <= 32'b10111100011000010110111011010100 ;
        3549: q <= 32'b10111100110000101000010001001111 ;
        3550: q <= 32'b00111101000110011100000101011100 ;
        3551: q <= 32'b00111101101000110000011110011101 ;
        3552: q <= 32'b00111101001001110101111000110001 ;
        3553: q <= 32'b10111011000010110110000110111111 ;
        3554: q <= 32'b00111100110111101010110010111000 ;
        3555: q <= 32'b00111101100101111111001110001000 ;
        3556: q <= 32'b10111101001100111001110110001101 ;
        3557: q <= 32'b00111100110010000010010100001000 ;
        3558: q <= 32'b00111100100111101101100101100001 ;
        3559: q <= 32'b10111100111010101110101100010110 ;
        3560: q <= 32'b00000000000000000000000000000000 ;
        3561: q <= 32'b00000000000000000000000000000000 ;
        3562: q <= 32'b00000000000000000000000000000000 ;
        3563: q <= 32'b00000000000000000000000000000000 ;
        3564: q <= 32'b00000000000000000000000000000000 ;
        3565: q <= 32'b00000000000000000000000000000000 ;
        3566: q <= 32'b00000000000000000000000000000000 ;
        3567: q <= 32'b00000000000000000000000000000000 ;
        3568: q <= 32'b00000000000000000000000000000000 ;
        3569: q <= 32'b00000000000000000000000000000000 ;
        3570: q <= 32'b00000000000000000000000000000000 ;
        3571: q <= 32'b00000000000000000000000000000000 ;
        3572: q <= 32'b00000000000000000000000000000000 ;
        3573: q <= 32'b00000000000000000000000000000000 ;
        3574: q <= 32'b00000000000000000000000000000000 ;
        3575: q <= 32'b00000000000000000000000000000000 ;
        3576: q <= 32'b00000000000000000000000000000000 ;
        3577: q <= 32'b00000000000000000000000000000000 ;
        3578: q <= 32'b00000000000000000000000000000000 ;
        3579: q <= 32'b00000000000000000000000000000000 ;
        3580: q <= 32'b00000000000000000000000000000000 ;
        3581: q <= 32'b00000000000000000000000000000000 ;
        3582: q <= 32'b00000000000000000000000000000000 ;
        3583: q <= 32'b00000000000000000000000000000000 ;
        3584: q <= 32'b00000000000000000000000000000000 ;
        3585: q <= 32'b00000000000000000000000000000000 ;
        3586: q <= 32'b00000000000000000000000000000000 ;
        3587: q <= 32'b00000000000000000000000000000000 ;
        3588: q <= 32'b00000000000000000000000000000000 ;
        3589: q <= 32'b00000000000000000000000000000000 ;
        3590: q <= 32'b00000000000000000000000000000000 ;
        3591: q <= 32'b00000000000000000000000000000000 ;
        3592: q <= 32'b00000000000000000000000000000000 ;
        3593: q <= 32'b00000000000000000000000000000000 ;
        3594: q <= 32'b00000000000000000000000000000000 ;
        3595: q <= 32'b00000000000000000000000000000000 ;
        3596: q <= 32'b00000000000000000000000000000000 ;
        3597: q <= 32'b00000000000000000000000000000000 ;
        3598: q <= 32'b00000000000000000000000000000000 ;
        3599: q <= 32'b00000000000000000000000000000000 ;
        3600: q <= 32'b00000000000000000000000000000000 ;
        3601: q <= 32'b00000000000000000000000000000000 ;
        3602: q <= 32'b00000000000000000000000000000000 ;
        3603: q <= 32'b00000000000000000000000000000000 ;
        3604: q <= 32'b00000000000000000000000000000000 ;
        3605: q <= 32'b00000000000000000000000000000000 ;
        3606: q <= 32'b00000000000000000000000000000000 ;
        3607: q <= 32'b00000000000000000000000000000000 ;
        3608: q <= 32'b00000000000000000000000000000000 ;
        3609: q <= 32'b00000000000000000000000000000000 ;
        3610: q <= 32'b00000000000000000000000000000000 ;
        3611: q <= 32'b00000000000000000000000000000000 ;
        3612: q <= 32'b00000000000000000000000000000000 ;
        3613: q <= 32'b00000000000000000000000000000000 ;
        3614: q <= 32'b00000000000000000000000000000000 ;
        3615: q <= 32'b00000000000000000000000000000000 ;
        3616: q <= 32'b00000000000000000000000000000000 ;
        3617: q <= 32'b00000000000000000000000000000000 ;
        3618: q <= 32'b00000000000000000000000000000000 ;
        3619: q <= 32'b00000000000000000000000000000000 ;
        3620: q <= 32'b00000000000000000000000000000000 ;
        3621: q <= 32'b00000000000000000000000000000000 ;
        3622: q <= 32'b00000000000000000000000000000000 ;
        3623: q <= 32'b00000000000000000000000000000000 ;
        3624: q <= 32'b00000000000000000000000000000000 ;
        3625: q <= 32'b00000000000000000000000000000000 ;
        3626: q <= 32'b00000000000000000000000000000000 ;
        3627: q <= 32'b00000000000000000000000000000000 ;
        3628: q <= 32'b00000000000000000000000000000000 ;
        3629: q <= 32'b00000000000000000000000000000000 ;
        3630: q <= 32'b00000000000000000000000000000000 ;
        3631: q <= 32'b00000000000000000000000000000000 ;
        3632: q <= 32'b00000000000000000000000000000000 ;
        3633: q <= 32'b00000000000000000000000000000000 ;
        3634: q <= 32'b00000000000000000000000000000000 ;
        3635: q <= 32'b00000000000000000000000000000000 ;
        3636: q <= 32'b00000000000000000000000000000000 ;
        3637: q <= 32'b00000000000000000000000000000000 ;
        3638: q <= 32'b00000000000000000000000000000000 ;
        3639: q <= 32'b00000000000000000000000000000000 ;
        3640: q <= 32'b00000000000000000000000000000000 ;
        3641: q <= 32'b00000000000000000000000000000000 ;
        3642: q <= 32'b00000000000000000000000000000000 ;
        3643: q <= 32'b00000000000000000000000000000000 ;
        3644: q <= 32'b00000000000000000000000000000000 ;
        3645: q <= 32'b00000000000000000000000000000000 ;
        3646: q <= 32'b00000000000000000000000000000000 ;
        3647: q <= 32'b00000000000000000000000000000000 ;
        3648: q <= 32'b00000000000000000000000000000000 ;
        3649: q <= 32'b00000000000000000000000000000000 ;
        3650: q <= 32'b00000000000000000000000000000000 ;
        3651: q <= 32'b00000000000000000000000000000000 ;
        3652: q <= 32'b00000000000000000000000000000000 ;
        3653: q <= 32'b00000000000000000000000000000000 ;
        3654: q <= 32'b00000000000000000000000000000000 ;
        3655: q <= 32'b00000000000000000000000000000000 ;
        3656: q <= 32'b00000000000000000000000000000000 ;
        3657: q <= 32'b00000000000000000000000000000000 ;
        3658: q <= 32'b00000000000000000000000000000000 ;
        3659: q <= 32'b00000000000000000000000000000000 ;
        3660: q <= 32'b00000000000000000000000000000000 ;
        3661: q <= 32'b00000000000000000000000000000000 ;
        3662: q <= 32'b00000000000000000000000000000000 ;
        3663: q <= 32'b00000000000000000000000000000000 ;
        3664: q <= 32'b00000000000000000000000000000000 ;
        3665: q <= 32'b00000000000000000000000000000000 ;
        3666: q <= 32'b00000000000000000000000000000000 ;
        3667: q <= 32'b00000000000000000000000000000000 ;
        3668: q <= 32'b00000000000000000000000000000000 ;
        3669: q <= 32'b00000000000000000000000000000000 ;
        3670: q <= 32'b00000000000000000000000000000000 ;
        3671: q <= 32'b00000000000000000000000000000000 ;
        3672: q <= 32'b00000000000000000000000000000000 ;
        3673: q <= 32'b00000000000000000000000000000000 ;
        3674: q <= 32'b00000000000000000000000000000000 ;
        3675: q <= 32'b00000000000000000000000000000000 ;
        3676: q <= 32'b00000000000000000000000000000000 ;
        3677: q <= 32'b00000000000000000000000000000000 ;
        3678: q <= 32'b00000000000000000000000000000000 ;
        3679: q <= 32'b00000000000000000000000000000000 ;
        3680: q <= 32'b00000000000000000000000000000000 ;
        3681: q <= 32'b00000000000000000000000000000000 ;
        3682: q <= 32'b00000000000000000000000000000000 ;
        3683: q <= 32'b00000000000000000000000000000000 ;
        3684: q <= 32'b00000000000000000000000000000000 ;
        3685: q <= 32'b00000000000000000000000000000000 ;
        3686: q <= 32'b00000000000000000000000000000000 ;
        3687: q <= 32'b00000000000000000000000000000000 ;
        3688: q <= 32'b00000000000000000000000000000000 ;
        3689: q <= 32'b00000000000000000000000000000000 ;
        3690: q <= 32'b00000000000000000000000000000000 ;
        3691: q <= 32'b00000000000000000000000000000000 ;
        3692: q <= 32'b00000000000000000000000000000000 ;
        3693: q <= 32'b00000000000000000000000000000000 ;
        3694: q <= 32'b00000000000000000000000000000000 ;
        3695: q <= 32'b00000000000000000000000000000000 ;
        3696: q <= 32'b00000000000000000000000000000000 ;
        3697: q <= 32'b00000000000000000000000000000000 ;
        3698: q <= 32'b00000000000000000000000000000000 ;
        3699: q <= 32'b00000000000000000000000000000000 ;
        3700: q <= 32'b00000000000000000000000000000000 ;
        3701: q <= 32'b00000000000000000000000000000000 ;
        3702: q <= 32'b00000000000000000000000000000000 ;
        3703: q <= 32'b00000000000000000000000000000000 ;
        3704: q <= 32'b00000000000000000000000000000000 ;
        3705: q <= 32'b00000000000000000000000000000000 ;
        3706: q <= 32'b00000000000000000000000000000000 ;
        3707: q <= 32'b00000000000000000000000000000000 ;
        3708: q <= 32'b00000000000000000000000000000000 ;
        3709: q <= 32'b00000000000000000000000000000000 ;
        3710: q <= 32'b00000000000000000000000000000000 ;
        3711: q <= 32'b00000000000000000000000000000000 ;
        3712: q <= 32'b00000000000000000000000000000000 ;
        3713: q <= 32'b00000000000000000000000000000000 ;
        3714: q <= 32'b00000000000000000000000000000000 ;
        3715: q <= 32'b00000000000000000000000000000000 ;
        3716: q <= 32'b00000000000000000000000000000000 ;
        3717: q <= 32'b00000000000000000000000000000000 ;
        3718: q <= 32'b00000000000000000000000000000000 ;
        3719: q <= 32'b00000000000000000000000000000000 ;
        3720: q <= 32'b00000000000000000000000000000000 ;
        3721: q <= 32'b00000000000000000000000000000000 ;
        3722: q <= 32'b00000000000000000000000000000000 ;
        3723: q <= 32'b00000000000000000000000000000000 ;
        3724: q <= 32'b00000000000000000000000000000000 ;
        3725: q <= 32'b00000000000000000000000000000000 ;
        3726: q <= 32'b00000000000000000000000000000000 ;
        3727: q <= 32'b00000000000000000000000000000000 ;
        3728: q <= 32'b00000000000000000000000000000000 ;
        3729: q <= 32'b00000000000000000000000000000000 ;
        3730: q <= 32'b00000000000000000000000000000000 ;
        3731: q <= 32'b00000000000000000000000000000000 ;
        3732: q <= 32'b00000000000000000000000000000000 ;
        3733: q <= 32'b00000000000000000000000000000000 ;
        3734: q <= 32'b00000000000000000000000000000000 ;
        3735: q <= 32'b00000000000000000000000000000000 ;
        3736: q <= 32'b00000000000000000000000000000000 ;
        3737: q <= 32'b00000000000000000000000000000000 ;
        3738: q <= 32'b00000000000000000000000000000000 ;
        3739: q <= 32'b00000000000000000000000000000000 ;
        3740: q <= 32'b00000000000000000000000000000000 ;
        3741: q <= 32'b00000000000000000000000000000000 ;
        3742: q <= 32'b00000000000000000000000000000000 ;
        3743: q <= 32'b00000000000000000000000000000000 ;
        3744: q <= 32'b00000000000000000000000000000000 ;
        3745: q <= 32'b00000000000000000000000000000000 ;
        3746: q <= 32'b00000000000000000000000000000000 ;
        3747: q <= 32'b00000000000000000000000000000000 ;
        3748: q <= 32'b00000000000000000000000000000000 ;
        3749: q <= 32'b00000000000000000000000000000000 ;
        3750: q <= 32'b00000000000000000000000000000000 ;
        3751: q <= 32'b00000000000000000000000000000000 ;
        3752: q <= 32'b00000000000000000000000000000000 ;
        3753: q <= 32'b00000000000000000000000000000000 ;
        3754: q <= 32'b00000000000000000000000000000000 ;
        3755: q <= 32'b00000000000000000000000000000000 ;
        3756: q <= 32'b00000000000000000000000000000000 ;
        3757: q <= 32'b00000000000000000000000000000000 ;
        3758: q <= 32'b00000000000000000000000000000000 ;
        3759: q <= 32'b00000000000000000000000000000000 ;
        3760: q <= 32'b00000000000000000000000000000000 ;
        3761: q <= 32'b00000000000000000000000000000000 ;
        3762: q <= 32'b00000000000000000000000000000000 ;
        3763: q <= 32'b00000000000000000000000000000000 ;
        3764: q <= 32'b00000000000000000000000000000000 ;
        3765: q <= 32'b00000000000000000000000000000000 ;
        3766: q <= 32'b00000000000000000000000000000000 ;
        3767: q <= 32'b00000000000000000000000000000000 ;
        3768: q <= 32'b00000000000000000000000000000000 ;
        3769: q <= 32'b00000000000000000000000000000000 ;
        3770: q <= 32'b00000000000000000000000000000000 ;
        3771: q <= 32'b00000000000000000000000000000000 ;
        3772: q <= 32'b00000000000000000000000000000000 ;
        3773: q <= 32'b00000000000000000000000000000000 ;
        3774: q <= 32'b00000000000000000000000000000000 ;
        3775: q <= 32'b00000000000000000000000000000000 ;
        3776: q <= 32'b00000000000000000000000000000000 ;
        3777: q <= 32'b00000000000000000000000000000000 ;
        3778: q <= 32'b00000000000000000000000000000000 ;
        3779: q <= 32'b00000000000000000000000000000000 ;
        3780: q <= 32'b00000000000000000000000000000000 ;
        3781: q <= 32'b00000000000000000000000000000000 ;
        3782: q <= 32'b00000000000000000000000000000000 ;
        3783: q <= 32'b00000000000000000000000000000000 ;
        3784: q <= 32'b00000000000000000000000000000000 ;
        3785: q <= 32'b00000000000000000000000000000000 ;
        3786: q <= 32'b00000000000000000000000000000000 ;
        3787: q <= 32'b00000000000000000000000000000000 ;
        3788: q <= 32'b00000000000000000000000000000000 ;
        3789: q <= 32'b00000000000000000000000000000000 ;
        3790: q <= 32'b00000000000000000000000000000000 ;
        3791: q <= 32'b00000000000000000000000000000000 ;
        3792: q <= 32'b00000000000000000000000000000000 ;
        3793: q <= 32'b00000000000000000000000000000000 ;
        3794: q <= 32'b00000000000000000000000000000000 ;
        3795: q <= 32'b00000000000000000000000000000000 ;
        3796: q <= 32'b00000000000000000000000000000000 ;
        3797: q <= 32'b00000000000000000000000000000000 ;
        3798: q <= 32'b00000000000000000000000000000000 ;
        3799: q <= 32'b00000000000000000000000000000000 ;
        3800: q <= 32'b00000000000000000000000000000000 ;
        3801: q <= 32'b00000000000000000000000000000000 ;
        3802: q <= 32'b00000000000000000000000000000000 ;
        3803: q <= 32'b00000000000000000000000000000000 ;
        3804: q <= 32'b00000000000000000000000000000000 ;
        3805: q <= 32'b00000000000000000000000000000000 ;
        3806: q <= 32'b00000000000000000000000000000000 ;
        3807: q <= 32'b00000000000000000000000000000000 ;
        3808: q <= 32'b00000000000000000000000000000000 ;
        3809: q <= 32'b00000000000000000000000000000000 ;
        3810: q <= 32'b00000000000000000000000000000000 ;
        3811: q <= 32'b00000000000000000000000000000000 ;
        3812: q <= 32'b00000000000000000000000000000000 ;
        3813: q <= 32'b00000000000000000000000000000000 ;
        3814: q <= 32'b00000000000000000000000000000000 ;
        3815: q <= 32'b00000000000000000000000000000000 ;
        3816: q <= 32'b00000000000000000000000000000000 ;
        3817: q <= 32'b00000000000000000000000000000000 ;
        3818: q <= 32'b00000000000000000000000000000000 ;
        3819: q <= 32'b00000000000000000000000000000000 ;
        3820: q <= 32'b00000000000000000000000000000000 ;
        3821: q <= 32'b00000000000000000000000000000000 ;
        3822: q <= 32'b00000000000000000000000000000000 ;
        3823: q <= 32'b00000000000000000000000000000000 ;
        3824: q <= 32'b00000000000000000000000000000000 ;
        3825: q <= 32'b00000000000000000000000000000000 ;
        3826: q <= 32'b00000000000000000000000000000000 ;
        3827: q <= 32'b00000000000000000000000000000000 ;
        3828: q <= 32'b00000000000000000000000000000000 ;
        3829: q <= 32'b00000000000000000000000000000000 ;
        3830: q <= 32'b00000000000000000000000000000000 ;
        3831: q <= 32'b00000000000000000000000000000000 ;
        3832: q <= 32'b00000000000000000000000000000000 ;
        3833: q <= 32'b00000000000000000000000000000000 ;
        3834: q <= 32'b00000000000000000000000000000000 ;
        3835: q <= 32'b00000000000000000000000000000000 ;
        3836: q <= 32'b00000000000000000000000000000000 ;
        3837: q <= 32'b00000000000000000000000000000000 ;
        3838: q <= 32'b00000000000000000000000000000000 ;
        3839: q <= 32'b00000000000000000000000000000000 ;
        3840: q <= 32'b00000000000000000000000000000000 ;
        3841: q <= 32'b00000000000000000000000000000000 ;
        3842: q <= 32'b00000000000000000000000000000000 ;
        3843: q <= 32'b00000000000000000000000000000000 ;
        3844: q <= 32'b00000000000000000000000000000000 ;
        3845: q <= 32'b00000000000000000000000000000000 ;
        3846: q <= 32'b00000000000000000000000000000000 ;
        3847: q <= 32'b00000000000000000000000000000000 ;
        3848: q <= 32'b00000000000000000000000000000000 ;
        3849: q <= 32'b00000000000000000000000000000000 ;
        3850: q <= 32'b00000000000000000000000000000000 ;
        3851: q <= 32'b00000000000000000000000000000000 ;
        3852: q <= 32'b00000000000000000000000000000000 ;
        3853: q <= 32'b00000000000000000000000000000000 ;
        3854: q <= 32'b00000000000000000000000000000000 ;
        3855: q <= 32'b00000000000000000000000000000000 ;
        3856: q <= 32'b00000000000000000000000000000000 ;
        3857: q <= 32'b00000000000000000000000000000000 ;
        3858: q <= 32'b00000000000000000000000000000000 ;
        3859: q <= 32'b00000000000000000000000000000000 ;
        3860: q <= 32'b00000000000000000000000000000000 ;
        3861: q <= 32'b00000000000000000000000000000000 ;
        3862: q <= 32'b00000000000000000000000000000000 ;
        3863: q <= 32'b00000000000000000000000000000000 ;
        3864: q <= 32'b00000000000000000000000000000000 ;
        3865: q <= 32'b00000000000000000000000000000000 ;
        3866: q <= 32'b00000000000000000000000000000000 ;
        3867: q <= 32'b00000000000000000000000000000000 ;
        3868: q <= 32'b00000000000000000000000000000000 ;
        3869: q <= 32'b00000000000000000000000000000000 ;
        3870: q <= 32'b00000000000000000000000000000000 ;
        3871: q <= 32'b00000000000000000000000000000000 ;
        3872: q <= 32'b00000000000000000000000000000000 ;
        3873: q <= 32'b00000000000000000000000000000000 ;
        3874: q <= 32'b00000000000000000000000000000000 ;
        3875: q <= 32'b00000000000000000000000000000000 ;
        3876: q <= 32'b00000000000000000000000000000000 ;
        3877: q <= 32'b00000000000000000000000000000000 ;
        3878: q <= 32'b00000000000000000000000000000000 ;
        3879: q <= 32'b00000000000000000000000000000000 ;
        3880: q <= 32'b00000000000000000000000000000000 ;
        3881: q <= 32'b00000000000000000000000000000000 ;
        3882: q <= 32'b00000000000000000000000000000000 ;
        3883: q <= 32'b00000000000000000000000000000000 ;
        3884: q <= 32'b00000000000000000000000000000000 ;
        3885: q <= 32'b00000000000000000000000000000000 ;
        3886: q <= 32'b00000000000000000000000000000000 ;
        3887: q <= 32'b00000000000000000000000000000000 ;
        3888: q <= 32'b00000000000000000000000000000000 ;
        3889: q <= 32'b00000000000000000000000000000000 ;
        3890: q <= 32'b00000000000000000000000000000000 ;
        3891: q <= 32'b00000000000000000000000000000000 ;
        3892: q <= 32'b00000000000000000000000000000000 ;
        3893: q <= 32'b00000000000000000000000000000000 ;
        3894: q <= 32'b00000000000000000000000000000000 ;
        3895: q <= 32'b00000000000000000000000000000000 ;
        3896: q <= 32'b00000000000000000000000000000000 ;
        3897: q <= 32'b00000000000000000000000000000000 ;
        3898: q <= 32'b00000000000000000000000000000000 ;
        3899: q <= 32'b00000000000000000000000000000000 ;
        3900: q <= 32'b00000000000000000000000000000000 ;
        3901: q <= 32'b00000000000000000000000000000000 ;
        3902: q <= 32'b00000000000000000000000000000000 ;
        3903: q <= 32'b00000000000000000000000000000000 ;
        3904: q <= 32'b00000000000000000000000000000000 ;
        3905: q <= 32'b00000000000000000000000000000000 ;
        3906: q <= 32'b00000000000000000000000000000000 ;
        3907: q <= 32'b00000000000000000000000000000000 ;
        3908: q <= 32'b00000000000000000000000000000000 ;
        3909: q <= 32'b00000000000000000000000000000000 ;
        3910: q <= 32'b00000000000000000000000000000000 ;
        3911: q <= 32'b00000000000000000000000000000000 ;
        3912: q <= 32'b00000000000000000000000000000000 ;
        3913: q <= 32'b00000000000000000000000000000000 ;
        3914: q <= 32'b00000000000000000000000000000000 ;
        3915: q <= 32'b00000000000000000000000000000000 ;
        3916: q <= 32'b00000000000000000000000000000000 ;
        3917: q <= 32'b00000000000000000000000000000000 ;
        3918: q <= 32'b00000000000000000000000000000000 ;
        3919: q <= 32'b00000000000000000000000000000000 ;
        3920: q <= 32'b00000000000000000000000000000000 ;
        3921: q <= 32'b00000000000000000000000000000000 ;
        3922: q <= 32'b00000000000000000000000000000000 ;
        3923: q <= 32'b00000000000000000000000000000000 ;
        3924: q <= 32'b00000000000000000000000000000000 ;
        3925: q <= 32'b00000000000000000000000000000000 ;
        3926: q <= 32'b00000000000000000000000000000000 ;
        3927: q <= 32'b00000000000000000000000000000000 ;
        3928: q <= 32'b00000000000000000000000000000000 ;
        3929: q <= 32'b00000000000000000000000000000000 ;
        3930: q <= 32'b00000000000000000000000000000000 ;
        3931: q <= 32'b00000000000000000000000000000000 ;
        3932: q <= 32'b00000000000000000000000000000000 ;
        3933: q <= 32'b00000000000000000000000000000000 ;
        3934: q <= 32'b00000000000000000000000000000000 ;
        3935: q <= 32'b00000000000000000000000000000000 ;
        3936: q <= 32'b00000000000000000000000000000000 ;
        3937: q <= 32'b00000000000000000000000000000000 ;
        3938: q <= 32'b00000000000000000000000000000000 ;
        3939: q <= 32'b00000000000000000000000000000000 ;
        3940: q <= 32'b00000000000000000000000000000000 ;
        3941: q <= 32'b00000000000000000000000000000000 ;
        3942: q <= 32'b00000000000000000000000000000000 ;
        3943: q <= 32'b00000000000000000000000000000000 ;
        3944: q <= 32'b00000000000000000000000000000000 ;
        3945: q <= 32'b00000000000000000000000000000000 ;
        3946: q <= 32'b00000000000000000000000000000000 ;
        3947: q <= 32'b00000000000000000000000000000000 ;
        3948: q <= 32'b00000000000000000000000000000000 ;
        3949: q <= 32'b00000000000000000000000000000000 ;
        3950: q <= 32'b00000000000000000000000000000000 ;
        3951: q <= 32'b00000000000000000000000000000000 ;
        3952: q <= 32'b00000000000000000000000000000000 ;
        3953: q <= 32'b00000000000000000000000000000000 ;
        3954: q <= 32'b00000000000000000000000000000000 ;
        3955: q <= 32'b00000000000000000000000000000000 ;
        3956: q <= 32'b00000000000000000000000000000000 ;
        3957: q <= 32'b00000000000000000000000000000000 ;
        3958: q <= 32'b00000000000000000000000000000000 ;
        3959: q <= 32'b00000000000000000000000000000000 ;
        3960: q <= 32'b00000000000000000000000000000000 ;
        3961: q <= 32'b00000000000000000000000000000000 ;
        3962: q <= 32'b00000000000000000000000000000000 ;
        3963: q <= 32'b00000000000000000000000000000000 ;
        3964: q <= 32'b00000000000000000000000000000000 ;
        3965: q <= 32'b00000000000000000000000000000000 ;
        3966: q <= 32'b00000000000000000000000000000000 ;
        3967: q <= 32'b00000000000000000000000000000000 ;
        3968: q <= 32'b00000000000000000000000000000000 ;
        3969: q <= 32'b00000000000000000000000000000000 ;
        3970: q <= 32'b00000000000000000000000000000000 ;
        3971: q <= 32'b00000000000000000000000000000000 ;
        3972: q <= 32'b00000000000000000000000000000000 ;
        3973: q <= 32'b00000000000000000000000000000000 ;
        3974: q <= 32'b00000000000000000000000000000000 ;
        3975: q <= 32'b00000000000000000000000000000000 ;
        3976: q <= 32'b00000000000000000000000000000000 ;
        3977: q <= 32'b00000000000000000000000000000000 ;
        3978: q <= 32'b00000000000000000000000000000000 ;
        3979: q <= 32'b00000000000000000000000000000000 ;
        3980: q <= 32'b00000000000000000000000000000000 ;
        3981: q <= 32'b00000000000000000000000000000000 ;
        3982: q <= 32'b00000000000000000000000000000000 ;
        3983: q <= 32'b00000000000000000000000000000000 ;
        3984: q <= 32'b00000000000000000000000000000000 ;
        3985: q <= 32'b00000000000000000000000000000000 ;
        3986: q <= 32'b00000000000000000000000000000000 ;
        3987: q <= 32'b00000000000000000000000000000000 ;
        3988: q <= 32'b00000000000000000000000000000000 ;
        3989: q <= 32'b00000000000000000000000000000000 ;
        3990: q <= 32'b00000000000000000000000000000000 ;
        3991: q <= 32'b00000000000000000000000000000000 ;
        3992: q <= 32'b00000000000000000000000000000000 ;
        3993: q <= 32'b00000000000000000000000000000000 ;
        3994: q <= 32'b00000000000000000000000000000000 ;
        3995: q <= 32'b00000000000000000000000000000000 ;
        3996: q <= 32'b00000000000000000000000000000000 ;
        3997: q <= 32'b00000000000000000000000000000000 ;
        3998: q <= 32'b00000000000000000000000000000000 ;
        3999: q <= 32'b00000000000000000000000000000000 ;
        4000: q <= 32'b00000000000000000000000000000000 ;
        4001: q <= 32'b00000000000000000000000000000000 ;
        4002: q <= 32'b00000000000000000000000000000000 ;
        4003: q <= 32'b00000000000000000000000000000000 ;
        4004: q <= 32'b00000000000000000000000000000000 ;
        4005: q <= 32'b00000000000000000000000000000000 ;
        4006: q <= 32'b00000000000000000000000000000000 ;
        4007: q <= 32'b00000000000000000000000000000000 ;
        4008: q <= 32'b00000000000000000000000000000000 ;
        4009: q <= 32'b00000000000000000000000000000000 ;
        4010: q <= 32'b00000000000000000000000000000000 ;
        4011: q <= 32'b00000000000000000000000000000000 ;
        4012: q <= 32'b00000000000000000000000000000000 ;
        4013: q <= 32'b00000000000000000000000000000000 ;
        4014: q <= 32'b00000000000000000000000000000000 ;
        4015: q <= 32'b00000000000000000000000000000000 ;
        4016: q <= 32'b00000000000000000000000000000000 ;
        4017: q <= 32'b00000000000000000000000000000000 ;
        4018: q <= 32'b00000000000000000000000000000000 ;
        4019: q <= 32'b00000000000000000000000000000000 ;
        4020: q <= 32'b00000000000000000000000000000000 ;
        4021: q <= 32'b00000000000000000000000000000000 ;
        4022: q <= 32'b00000000000000000000000000000000 ;
        4023: q <= 32'b00000000000000000000000000000000 ;
        4024: q <= 32'b00000000000000000000000000000000 ;
        4025: q <= 32'b00000000000000000000000000000000 ;
        4026: q <= 32'b00000000000000000000000000000000 ;
        4027: q <= 32'b00000000000000000000000000000000 ;
        4028: q <= 32'b00000000000000000000000000000000 ;
        4029: q <= 32'b00000000000000000000000000000000 ;
        4030: q <= 32'b00000000000000000000000000000000 ;
        4031: q <= 32'b00000000000000000000000000000000 ;
        4032: q <= 32'b00000000000000000000000000000000 ;
        4033: q <= 32'b00000000000000000000000000000000 ;
        4034: q <= 32'b00000000000000000000000000000000 ;
        4035: q <= 32'b00000000000000000000000000000000 ;
        4036: q <= 32'b00000000000000000000000000000000 ;
        4037: q <= 32'b00000000000000000000000000000000 ;
        4038: q <= 32'b00000000000000000000000000000000 ;
        4039: q <= 32'b00000000000000000000000000000000 ;
        4040: q <= 32'b00000000000000000000000000000000 ;
        4041: q <= 32'b00000000000000000000000000000000 ;
        4042: q <= 32'b00000000000000000000000000000000 ;
        4043: q <= 32'b00000000000000000000000000000000 ;
        4044: q <= 32'b00000000000000000000000000000000 ;
        4045: q <= 32'b00000000000000000000000000000000 ;
        4046: q <= 32'b00000000000000000000000000000000 ;
        4047: q <= 32'b00000000000000000000000000000000 ;
        4048: q <= 32'b00000000000000000000000000000000 ;
        4049: q <= 32'b00000000000000000000000000000000 ;
        4050: q <= 32'b00000000000000000000000000000000 ;
        4051: q <= 32'b00000000000000000000000000000000 ;
        4052: q <= 32'b00000000000000000000000000000000 ;
        4053: q <= 32'b00000000000000000000000000000000 ;
        4054: q <= 32'b00000000000000000000000000000000 ;
        4055: q <= 32'b00000000000000000000000000000000 ;
        4056: q <= 32'b00000000000000000000000000000000 ;
        4057: q <= 32'b00000000000000000000000000000000 ;
        4058: q <= 32'b00000000000000000000000000000000 ;
        4059: q <= 32'b00000000000000000000000000000000 ;
        4060: q <= 32'b00000000000000000000000000000000 ;
        4061: q <= 32'b00000000000000000000000000000000 ;
        4062: q <= 32'b00000000000000000000000000000000 ;
        4063: q <= 32'b00000000000000000000000000000000 ;
        4064: q <= 32'b00000000000000000000000000000000 ;
        4065: q <= 32'b00000000000000000000000000000000 ;
        4066: q <= 32'b00000000000000000000000000000000 ;
        4067: q <= 32'b00000000000000000000000000000000 ;
        4068: q <= 32'b00000000000000000000000000000000 ;
        4069: q <= 32'b00000000000000000000000000000000 ;
        4070: q <= 32'b00000000000000000000000000000000 ;
        4071: q <= 32'b00000000000000000000000000000000 ;
        4072: q <= 32'b00000000000000000000000000000000 ;
        4073: q <= 32'b00000000000000000000000000000000 ;
        4074: q <= 32'b00000000000000000000000000000000 ;
        4075: q <= 32'b00000000000000000000000000000000 ;
        4076: q <= 32'b00000000000000000000000000000000 ;
        4077: q <= 32'b00000000000000000000000000000000 ;
        4078: q <= 32'b00000000000000000000000000000000 ;
        4079: q <= 32'b00000000000000000000000000000000 ;
        4080: q <= 32'b00000000000000000000000000000000 ;
        4081: q <= 32'b00000000000000000000000000000000 ;
        4082: q <= 32'b00000000000000000000000000000000 ;
        4083: q <= 32'b00000000000000000000000000000000 ;
        4084: q <= 32'b00000000000000000000000000000000 ;
        4085: q <= 32'b00000000000000000000000000000000 ;
        4086: q <= 32'b00000000000000000000000000000000 ;
        4087: q <= 32'b00000000000000000000000000000000 ;
        4088: q <= 32'b00000000000000000000000000000000 ;
        4089: q <= 32'b00000000000000000000000000000000 ;
        4090: q <= 32'b00000000000000000000000000000000 ;
        4091: q <= 32'b00000000000000000000000000000000 ;
        4092: q <= 32'b00000000000000000000000000000000 ;
        4093: q <= 32'b00000000000000000000000000000000 ;
        4094: q <= 32'b00000000000000000000000000000000 ;
        4095: q <= 32'b00000000000000000000000000000000 ;
        default: q <= 32'b00000000000000000000000000000000;
    endcase
end

endmodule
