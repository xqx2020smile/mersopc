module mem_rom_weight_out (clock, address, q) ;
parameter DATA_WIDTH =  32;
input clock;
input [10:0] address;
output [DATA_WIDTH-1:0] q;
reg    [DATA_WIDTH-1:0] q;
always@(posedge clock) begin 
    case(address)
        0: q <= 32'b00111101110000111000101110000001 ;
        1: q <= 32'b00111110001000011010001010001010 ;
        2: q <= 32'b10111110100010110110100111001001 ;
        3: q <= 32'b00111101110000001110000001101010 ;
        4: q <= 32'b00111110000111110001101100010000 ;
        5: q <= 32'b10111101110111110101011000101001 ;
        6: q <= 32'b10111110101010000110111100110001 ;
        7: q <= 32'b10111110100110110101110001110111 ;
        8: q <= 32'b00111101111010111110111110111010 ;
        9: q <= 32'b10111110100001011010100101001101 ;
        10: q <= 32'b10111111011100110100000000111001 ;
        11: q <= 32'b00111110010000000111100110101110 ;
        12: q <= 32'b10111110100100111011011001110011 ;
        13: q <= 32'b10111110100011000001101001100011 ;
        14: q <= 32'b10111111010011011101110101001111 ;
        15: q <= 32'b00111101100001111001111000111001 ;
        16: q <= 32'b10111110101110001001010001110010 ;
        17: q <= 32'b00111110010000100111111011110000 ;
        18: q <= 32'b10111111010010100001001101110000 ;
        19: q <= 32'b00111101001001100101100110100010 ;
        20: q <= 32'b10111111001011101100100011110111 ;
        21: q <= 32'b00111110110111000011001100011110 ;
        22: q <= 32'b10111110010011100011000010100010 ;
        23: q <= 32'b00111101110011111101000111100001 ;
        24: q <= 32'b10111110011110110111000011101010 ;
        25: q <= 32'b10111110001000100000100000110010 ;
        26: q <= 32'b10111110101110100110101100001001 ;
        27: q <= 32'b00111110100101111011101111000010 ;
        28: q <= 32'b10111110000111111110110001101011 ;
        29: q <= 32'b10111110100011010001111110110010 ;
        30: q <= 32'b00111101011101100101111101010000 ;
        31: q <= 32'b10111101111101010011101101110100 ;
        32: q <= 32'b10111110110110100011001011000110 ;
        33: q <= 32'b10111111010010100001000010000001 ;
        34: q <= 32'b00111111001110110110010001111010 ;
        35: q <= 32'b10111101001001011100000010110000 ;
        36: q <= 32'b00111110001111101001000110001111 ;
        37: q <= 32'b00111110101110000111100111101111 ;
        38: q <= 32'b00111011101000100010110111111011 ;
        39: q <= 32'b00111111000010100001011010100100 ;
        40: q <= 32'b00111100010001011001101101101100 ;
        41: q <= 32'b10111110101000111100110110110100 ;
        42: q <= 32'b00111110000000101111111010010101 ;
        43: q <= 32'b00111110000000101000100000111010 ;
        44: q <= 32'b10111110010000101010011011011010 ;
        45: q <= 32'b10111111001100111000111001110001 ;
        46: q <= 32'b10111110000101010011101010011010 ;
        47: q <= 32'b10111101100101100100110100100111 ;
        48: q <= 32'b00111110110010100101010011001000 ;
        49: q <= 32'b10111101111010110110000010000101 ;
        50: q <= 32'b10111110011100010001001111000001 ;
        51: q <= 32'b10111110101111110000101111100011 ;
        52: q <= 32'b00111110001110100110110001000111 ;
        53: q <= 32'b10111110111011000001100110000101 ;
        54: q <= 32'b10111101001000011010110100101010 ;
        55: q <= 32'b00111111001111001111001101111000 ;
        56: q <= 32'b00111110001101001010010100010000 ;
        57: q <= 32'b10111101000000001000101110010100 ;
        58: q <= 32'b00111110011001101001010000000111 ;
        59: q <= 32'b10111110100110010100111010011100 ;
        60: q <= 32'b00000000000000000000000000000000 ;
        61: q <= 32'b00000000000000000000000000000000 ;
        62: q <= 32'b00000000000000000000000000000000 ;
        63: q <= 32'b00000000000000000000000000000000 ;
        64: q <= 32'b10111110000011101110110111000011 ;
        65: q <= 32'b10111101000011111001000011010001 ;
        66: q <= 32'b10111011000000110110111011111100 ;
        67: q <= 32'b10111111001101011001011111010011 ;
        68: q <= 32'b00111101111000010111111011010000 ;
        69: q <= 32'b10111101100010000100000010111001 ;
        70: q <= 32'b00111110000011010011001000100100 ;
        71: q <= 32'b10111110011111000001100001110010 ;
        72: q <= 32'b00111101000111000000110001110011 ;
        73: q <= 32'b10111110100011111110101101111111 ;
        74: q <= 32'b10111110111011010011101110110100 ;
        75: q <= 32'b10111111001110100110011100001110 ;
        76: q <= 32'b00111110001100001011100101011111 ;
        77: q <= 32'b10111110010000010000110100001000 ;
        78: q <= 32'b10111111000010111000001001100111 ;
        79: q <= 32'b00111101101000001111110100111101 ;
        80: q <= 32'b10111110101111101010001000111000 ;
        81: q <= 32'b00111110001000101010011011101111 ;
        82: q <= 32'b00111110110001011000111110010001 ;
        83: q <= 32'b00111101111000010011001111011100 ;
        84: q <= 32'b00111110101010000110111101001101 ;
        85: q <= 32'b00111110001100101011000111101001 ;
        86: q <= 32'b00111111000110011011100111101100 ;
        87: q <= 32'b00111101110110101110011000010101 ;
        88: q <= 32'b10111110100010110010010011111010 ;
        89: q <= 32'b00111101011011000010000100011110 ;
        90: q <= 32'b00111111000000101100001010000000 ;
        91: q <= 32'b00111110001011110111101010001011 ;
        92: q <= 32'b00111110000100100011010001011111 ;
        93: q <= 32'b10111110010110000111111111100111 ;
        94: q <= 32'b00111110011100101001011111000001 ;
        95: q <= 32'b10111110000001010001111010110001 ;
        96: q <= 32'b10111110010110001011111100101110 ;
        97: q <= 32'b10111011011111010111100110001010 ;
        98: q <= 32'b00111110101101101011011100011101 ;
        99: q <= 32'b10111101110111000000111001101000 ;
        100: q <= 32'b10111101111111110010011010100101 ;
        101: q <= 32'b10111101101101001011000101001111 ;
        102: q <= 32'b10111111001000000000010101001000 ;
        103: q <= 32'b10111101111011011000111101100001 ;
        104: q <= 32'b10111100100000111110001101111100 ;
        105: q <= 32'b00111110010001000011101000000111 ;
        106: q <= 32'b00111110001010111110001001111100 ;
        107: q <= 32'b10111110111110000010100100010011 ;
        108: q <= 32'b10111110010011011101100100100101 ;
        109: q <= 32'b10111111001001101001101110100000 ;
        110: q <= 32'b10111110011010100000111111110011 ;
        111: q <= 32'b10111101011010010110011111001111 ;
        112: q <= 32'b10111110111011101011110100001110 ;
        113: q <= 32'b10111101111011111001111101101111 ;
        114: q <= 32'b10111101110111010000111010000100 ;
        115: q <= 32'b10111101011111100101011000101010 ;
        116: q <= 32'b00111110001010110000001011001110 ;
        117: q <= 32'b10111110011101101101110111110111 ;
        118: q <= 32'b00111100101011100010111111000011 ;
        119: q <= 32'b10111110010100000101001001000111 ;
        120: q <= 32'b00111110100100001101111000100110 ;
        121: q <= 32'b00111110010010100011001000000101 ;
        122: q <= 32'b00111110011101000011000011011110 ;
        123: q <= 32'b10111110011000110011110100111110 ;
        124: q <= 32'b00000000000000000000000000000000 ;
        125: q <= 32'b00000000000000000000000000000000 ;
        126: q <= 32'b00000000000000000000000000000000 ;
        127: q <= 32'b00000000000000000000000000000000 ;
        128: q <= 32'b10111101100001111010001111110011 ;
        129: q <= 32'b10111111000100011001000011101111 ;
        130: q <= 32'b00111110000110000110001110100110 ;
        131: q <= 32'b10111110000000000001001100100000 ;
        132: q <= 32'b00111110010000110100001111010010 ;
        133: q <= 32'b10111110001110001000101110101010 ;
        134: q <= 32'b00111010100011001101100011110110 ;
        135: q <= 32'b10111110101010000011011010001100 ;
        136: q <= 32'b10111101101010001100100000000001 ;
        137: q <= 32'b10111101111000101001011011011001 ;
        138: q <= 32'b00111110001110010101100100011110 ;
        139: q <= 32'b10111101110100010100011111101001 ;
        140: q <= 32'b10111111001000001100101101101101 ;
        141: q <= 32'b10111110011011111100011011001110 ;
        142: q <= 32'b00111110001011010010110001100001 ;
        143: q <= 32'b00111110100111111101000011010111 ;
        144: q <= 32'b00111110101011101101111101111010 ;
        145: q <= 32'b00111110100001100111011010000010 ;
        146: q <= 32'b10111110101100011000010000110000 ;
        147: q <= 32'b00111110011111100110011101100100 ;
        148: q <= 32'b10111110101000111110110111100011 ;
        149: q <= 32'b00111110100010101100010000111110 ;
        150: q <= 32'b00111111001010110101010100101110 ;
        151: q <= 32'b00111101101011110000001011101111 ;
        152: q <= 32'b10111111001110100101101010111000 ;
        153: q <= 32'b10111100100011110100110111111011 ;
        154: q <= 32'b00111111000111111100110111000101 ;
        155: q <= 32'b00111110100101001110010001010000 ;
        156: q <= 32'b00111111001011000000101000001011 ;
        157: q <= 32'b10111110000001101101001001011001 ;
        158: q <= 32'b00111111010101001001001010001110 ;
        159: q <= 32'b10111110101001010000111001001010 ;
        160: q <= 32'b00111110011000111100001100110101 ;
        161: q <= 32'b00111101001101100111100000100011 ;
        162: q <= 32'b00111111001001101100100000101101 ;
        163: q <= 32'b10111111010000000011101101010101 ;
        164: q <= 32'b00111101110010101111100111010000 ;
        165: q <= 32'b00111100011000100111111001110001 ;
        166: q <= 32'b00111101100110100010101101001000 ;
        167: q <= 32'b00111110111111001110100100010010 ;
        168: q <= 32'b10111110000010100100111011000001 ;
        169: q <= 32'b10111111000011110010101101111001 ;
        170: q <= 32'b00111110001010010011011000010000 ;
        171: q <= 32'b00111101100000000010010000110110 ;
        172: q <= 32'b10111110000010111011101011010000 ;
        173: q <= 32'b00111101100001001011000011101000 ;
        174: q <= 32'b10111110011000011100111110101010 ;
        175: q <= 32'b00111101100001100000110000010000 ;
        176: q <= 32'b00111110001011101110111101010001 ;
        177: q <= 32'b10111110100000101000000011011100 ;
        178: q <= 32'b10111110100010101100111111000100 ;
        179: q <= 32'b00111111001001101000101011010111 ;
        180: q <= 32'b00111110001110111000011000100010 ;
        181: q <= 32'b10111101110110000100110101111101 ;
        182: q <= 32'b00111110011010101011010111110000 ;
        183: q <= 32'b10111110000001110100101000011100 ;
        184: q <= 32'b00111110101011011000000010100101 ;
        185: q <= 32'b10111101110001010111111010101100 ;
        186: q <= 32'b00111110100010100101101011011000 ;
        187: q <= 32'b10111101111000000001010111101010 ;
        188: q <= 32'b00000000000000000000000000000000 ;
        189: q <= 32'b00000000000000000000000000000000 ;
        190: q <= 32'b00000000000000000000000000000000 ;
        191: q <= 32'b00000000000000000000000000000000 ;
        192: q <= 32'b00111111000110011101000000000100 ;
        193: q <= 32'b00111101011110010011011001110110 ;
        194: q <= 32'b10111100111101010001000001011000 ;
        195: q <= 32'b00111101100000100001100101000000 ;
        196: q <= 32'b10111101001001011111100010110100 ;
        197: q <= 32'b10111110001100100001000101011101 ;
        198: q <= 32'b10111101110100100000111010000001 ;
        199: q <= 32'b10111110100000000010110110111110 ;
        200: q <= 32'b00111111010100110001000011000010 ;
        201: q <= 32'b10111101110100001010011110011010 ;
        202: q <= 32'b10111111001101101000001011001110 ;
        203: q <= 32'b00111101110100011001000001110110 ;
        204: q <= 32'b00111110101001110110010001101111 ;
        205: q <= 32'b10111110011000100101100110111110 ;
        206: q <= 32'b00111110100110100110001111101000 ;
        207: q <= 32'b00111110001000010010111000001011 ;
        208: q <= 32'b00111110101110111010100010110110 ;
        209: q <= 32'b00111101010010100100010101010011 ;
        210: q <= 32'b00111110100010111011011100011100 ;
        211: q <= 32'b00111110100100001001000010110001 ;
        212: q <= 32'b00111111000101110111001011111111 ;
        213: q <= 32'b00111110100110100000111011111110 ;
        214: q <= 32'b00111100100101011000010100101101 ;
        215: q <= 32'b00111111010111011110011101001110 ;
        216: q <= 32'b00111110100110000101100010001110 ;
        217: q <= 32'b00111100001110000110101011011000 ;
        218: q <= 32'b10111110010110100111000000011010 ;
        219: q <= 32'b00111101111010011111000010011100 ;
        220: q <= 32'b10111110000010001010011001100010 ;
        221: q <= 32'b10111101111010101110001100000000 ;
        222: q <= 32'b00111101100011100111001001100011 ;
        223: q <= 32'b10111111000110111111011101101011 ;
        224: q <= 32'b10111110100101011010100100101001 ;
        225: q <= 32'b10111100100100101111011000100011 ;
        226: q <= 32'b10111110100001101110010001111111 ;
        227: q <= 32'b10111101011001001111011101101000 ;
        228: q <= 32'b00111110011110011001011110010111 ;
        229: q <= 32'b00111110010110000101001101011110 ;
        230: q <= 32'b10111101001100000011000110010010 ;
        231: q <= 32'b00111111000110111100110011010010 ;
        232: q <= 32'b10111110001011000101100100101100 ;
        233: q <= 32'b00111101110000110010111010011011 ;
        234: q <= 32'b00111110000010110010010100010010 ;
        235: q <= 32'b10111110110110000110111011011000 ;
        236: q <= 32'b10111110100000010001111000111110 ;
        237: q <= 32'b10111101011010001011111111010010 ;
        238: q <= 32'b10111110011100001000111101111010 ;
        239: q <= 32'b10111101101101000001111111100001 ;
        240: q <= 32'b10111111001111101011100100011001 ;
        241: q <= 32'b10111101110101011101011110100101 ;
        242: q <= 32'b10111110101011010001000010100000 ;
        243: q <= 32'b00111101100111101010010010000010 ;
        244: q <= 32'b00111110010110010010001111110111 ;
        245: q <= 32'b10111101111000111010001111001101 ;
        246: q <= 32'b00111110001100000110000001100110 ;
        247: q <= 32'b00111110001110100001110101101101 ;
        248: q <= 32'b00111101111111111011111011101111 ;
        249: q <= 32'b10111101011000111110011011011110 ;
        250: q <= 32'b00111110100100111011110001001111 ;
        251: q <= 32'b10111110100000100011110100010111 ;
        252: q <= 32'b00000000000000000000000000000000 ;
        253: q <= 32'b00000000000000000000000000000000 ;
        254: q <= 32'b00000000000000000000000000000000 ;
        255: q <= 32'b00000000000000000000000000000000 ;
        256: q <= 32'b00111101111010101110000101111111 ;
        257: q <= 32'b10111101001110011000011110111010 ;
        258: q <= 32'b10111110000001010101101001011000 ;
        259: q <= 32'b00111101101100011000011100011011 ;
        260: q <= 32'b00111110001011101110010101100011 ;
        261: q <= 32'b10111101110011100000111000011111 ;
        262: q <= 32'b00111101110011110000100111000010 ;
        263: q <= 32'b10111110000111111001011111011010 ;
        264: q <= 32'b10111101010100110010011000110111 ;
        265: q <= 32'b10111110010000000111001011011101 ;
        266: q <= 32'b10111110111101110010011101111110 ;
        267: q <= 32'b10111111000000111110101011101101 ;
        268: q <= 32'b00111110011001111001111101101011 ;
        269: q <= 32'b10111110010011110111000010110000 ;
        270: q <= 32'b00111101111100010001110011000111 ;
        271: q <= 32'b00111101110000000001110000001010 ;
        272: q <= 32'b10111111000011111101101110010010 ;
        273: q <= 32'b10111100101000001001100000011101 ;
        274: q <= 32'b10111110101110010011010111000110 ;
        275: q <= 32'b00111110010101110110101111101011 ;
        276: q <= 32'b00111110110000111001110111000110 ;
        277: q <= 32'b00111110011001000000100101111101 ;
        278: q <= 32'b10111110001001101101111010111010 ;
        279: q <= 32'b00111110000110101101110001001011 ;
        280: q <= 32'b00111101110100010111001001110010 ;
        281: q <= 32'b10111110101100000111111000010111 ;
        282: q <= 32'b00111110110110001100111001011101 ;
        283: q <= 32'b00111110010000101101110000011110 ;
        284: q <= 32'b00111101101011100011001111001001 ;
        285: q <= 32'b10111110000001011100101011100111 ;
        286: q <= 32'b00111110100000111001101101101010 ;
        287: q <= 32'b10111101011011010011101101100111 ;
        288: q <= 32'b00111111000011000100100001110111 ;
        289: q <= 32'b10111100110100101110100000011100 ;
        290: q <= 32'b00111110101111010000010001010110 ;
        291: q <= 32'b10111110000010001011100101010011 ;
        292: q <= 32'b00111111010111001001010001100111 ;
        293: q <= 32'b00111111000101000100011101000011 ;
        294: q <= 32'b00111101101110101111101011011000 ;
        295: q <= 32'b10111110001011101100000111111000 ;
        296: q <= 32'b10111101001110100111011100010111 ;
        297: q <= 32'b10111110010111011001111110011111 ;
        298: q <= 32'b10111100110101000000000100111001 ;
        299: q <= 32'b00111110100111111100011101011001 ;
        300: q <= 32'b10111110100100111000001001101111 ;
        301: q <= 32'b00111110010000001000110010111000 ;
        302: q <= 32'b10111011100101010010010111101010 ;
        303: q <= 32'b10111101101100011111111001000001 ;
        304: q <= 32'b10111111000001110011001001000010 ;
        305: q <= 32'b10111110001100100110110000101101 ;
        306: q <= 32'b10111110100000100101010110101011 ;
        307: q <= 32'b00111110110100101010000000011100 ;
        308: q <= 32'b10111100101111101001010011010010 ;
        309: q <= 32'b00111111000110000111000010100000 ;
        310: q <= 32'b00111101101001100111100101110010 ;
        311: q <= 32'b00111110110000100110110010011001 ;
        312: q <= 32'b00111110010010011001001010000100 ;
        313: q <= 32'b10111111000001010111011101001001 ;
        314: q <= 32'b00111110001011111100011000010101 ;
        315: q <= 32'b10111101110111000000111001100000 ;
        316: q <= 32'b00000000000000000000000000000000 ;
        317: q <= 32'b00000000000000000000000000000000 ;
        318: q <= 32'b00000000000000000000000000000000 ;
        319: q <= 32'b00000000000000000000000000000000 ;
        320: q <= 32'b00111111010011101110001110011110 ;
        321: q <= 32'b10111111001011000010111101010111 ;
        322: q <= 32'b10111101100100001101100110110001 ;
        323: q <= 32'b10111101100100100011001110010000 ;
        324: q <= 32'b00111110001111010011011001011111 ;
        325: q <= 32'b10111110000100111000110011101011 ;
        326: q <= 32'b00111101001100110110110101101000 ;
        327: q <= 32'b10111110101100010100101101010100 ;
        328: q <= 32'b10111110001000010001000010001001 ;
        329: q <= 32'b10111110100000001010011101000111 ;
        330: q <= 32'b00111101100010110101011001001010 ;
        331: q <= 32'b10111101101100101000100100110111 ;
        332: q <= 32'b00111110111000111011110111100010 ;
        333: q <= 32'b10111110001010001000101100100101 ;
        334: q <= 32'b10111111010011111010111101011001 ;
        335: q <= 32'b00111110010111101101010000100010 ;
        336: q <= 32'b00111110000111011110011111010111 ;
        337: q <= 32'b00111101001001000011110010010110 ;
        338: q <= 32'b00111110111111111000100000000001 ;
        339: q <= 32'b00111110110100101100111100010101 ;
        340: q <= 32'b10111111000111000101011010110011 ;
        341: q <= 32'b00111110100100111010000101111110 ;
        342: q <= 32'b10111101101000001110111001000011 ;
        343: q <= 32'b00111100111001111000100101010110 ;
        344: q <= 32'b10111110111010111010010010101001 ;
        345: q <= 32'b00111100101001010011001110101101 ;
        346: q <= 32'b10111110110001101010111001011001 ;
        347: q <= 32'b00111110001100111101100111101000 ;
        348: q <= 32'b00111111001001001101111101001101 ;
        349: q <= 32'b10111101011100010110011110010111 ;
        350: q <= 32'b00111101010110000011110111110001 ;
        351: q <= 32'b00111110101010010101011000111100 ;
        352: q <= 32'b10111110100010011010001011111001 ;
        353: q <= 32'b10111110001111101000100000011010 ;
        354: q <= 32'b10111110101011010110010010000110 ;
        355: q <= 32'b10111111011100000000111111100100 ;
        356: q <= 32'b00111110101010010100011011111001 ;
        357: q <= 32'b10111101001101101101111101000101 ;
        358: q <= 32'b10111110010101111101001110010101 ;
        359: q <= 32'b00111111001000000101101101110100 ;
        360: q <= 32'b10111101100111111111100111111001 ;
        361: q <= 32'b00111110101000011001010100100111 ;
        362: q <= 32'b00111100100010010101011011000011 ;
        363: q <= 32'b10111111010011100001011010000111 ;
        364: q <= 32'b10111110011010010001000010101111 ;
        365: q <= 32'b00111101110101001001000111010111 ;
        366: q <= 32'b10111110101011110001101111011011 ;
        367: q <= 32'b10111110001001001110001111100110 ;
        368: q <= 32'b00111110001000010011000000001000 ;
        369: q <= 32'b10111110000101110100101010101010 ;
        370: q <= 32'b10111110101001001110001001101011 ;
        371: q <= 32'b00111101111011010011100100100101 ;
        372: q <= 32'b00111110010011101011111001011101 ;
        373: q <= 32'b00111101110101010010111000101111 ;
        374: q <= 32'b00111110001010111101000100000010 ;
        375: q <= 32'b00111110010110011011100100101011 ;
        376: q <= 32'b00111110001001000000110011000111 ;
        377: q <= 32'b00111101010101001010011110100010 ;
        378: q <= 32'b00111110101101100000111010000000 ;
        379: q <= 32'b10111110001111011010000100101011 ;
        380: q <= 32'b00000000000000000000000000000000 ;
        381: q <= 32'b00000000000000000000000000000000 ;
        382: q <= 32'b00000000000000000000000000000000 ;
        383: q <= 32'b00000000000000000000000000000000 ;
        384: q <= 32'b00111111000100111010101111100001 ;
        385: q <= 32'b10111110000001001100000010111110 ;
        386: q <= 32'b10111110101001010101101001110111 ;
        387: q <= 32'b00111110000100011111100101110000 ;
        388: q <= 32'b00111111011100010010111000010100 ;
        389: q <= 32'b10111110100000000000000011100010 ;
        390: q <= 32'b00111101101101010001111100100011 ;
        391: q <= 32'b10111110001010010110101010111010 ;
        392: q <= 32'b10111101100001011111011110111011 ;
        393: q <= 32'b10111110001001110110011110011010 ;
        394: q <= 32'b00111110101000011001111110111110 ;
        395: q <= 32'b00111110001010100001101010001001 ;
        396: q <= 32'b00111110010000010010101010101110 ;
        397: q <= 32'b10111110100001110000001111001011 ;
        398: q <= 32'b00111110101011101111110101100110 ;
        399: q <= 32'b00111110010000110100100011110111 ;
        400: q <= 32'b00111110011010111111000110110100 ;
        401: q <= 32'b00111101110100110111101101111100 ;
        402: q <= 32'b10111110111111000110001100000001 ;
        403: q <= 32'b00111110011011011111100010110011 ;
        404: q <= 32'b00111101011011001011111111110111 ;
        405: q <= 32'b00111101000000101011101000001100 ;
        406: q <= 32'b00111011100010100000011001010111 ;
        407: q <= 32'b00111100101100110000011100110001 ;
        408: q <= 32'b10111110111000101010001111011001 ;
        409: q <= 32'b10111110000011010100111111101000 ;
        410: q <= 32'b10111110111001010100000000001011 ;
        411: q <= 32'b00111110100011101001010101101111 ;
        412: q <= 32'b10111110011001000011111100100000 ;
        413: q <= 32'b10111110010101110100111101010110 ;
        414: q <= 32'b00111101101011011101001100001011 ;
        415: q <= 32'b00111110101100001101111100111110 ;
        416: q <= 32'b10111101111110010111010110100001 ;
        417: q <= 32'b10111100110100111110101010111111 ;
        418: q <= 32'b00111111000000101110100001001000 ;
        419: q <= 32'b10111101100000111100100110010111 ;
        420: q <= 32'b00111100110011111000010010101000 ;
        421: q <= 32'b10111110011001000000101101010101 ;
        422: q <= 32'b00111110000100110110111100110101 ;
        423: q <= 32'b10111110110001010111101101011100 ;
        424: q <= 32'b10111111001110101011101000110000 ;
        425: q <= 32'b00111110100110111010100010110111 ;
        426: q <= 32'b00111110010111001000010010111000 ;
        427: q <= 32'b00111110111100000100101111111011 ;
        428: q <= 32'b10111110100010000100011101010111 ;
        429: q <= 32'b10111111010111010000110010111010 ;
        430: q <= 32'b10111110000111100011011100011101 ;
        431: q <= 32'b10111101001110010000000111111111 ;
        432: q <= 32'b10111111001101101001010101111011 ;
        433: q <= 32'b10111110000111110001001001011111 ;
        434: q <= 32'b10111110000010000000000010000011 ;
        435: q <= 32'b00111111010100000000010001010110 ;
        436: q <= 32'b00111110011100101001001100001110 ;
        437: q <= 32'b00111101100110100100001100111000 ;
        438: q <= 32'b10111111001001010100101001001110 ;
        439: q <= 32'b10111110000001110100100001011110 ;
        440: q <= 32'b00111110010001010000010010100001 ;
        441: q <= 32'b00111100101101010011011100110011 ;
        442: q <= 32'b00111110100000111110010111110111 ;
        443: q <= 32'b10111110010101001000110001010100 ;
        444: q <= 32'b00000000000000000000000000000000 ;
        445: q <= 32'b00000000000000000000000000000000 ;
        446: q <= 32'b00000000000000000000000000000000 ;
        447: q <= 32'b00000000000000000000000000000000 ;
        448: q <= 32'b00111100110011001101101100000000 ;
        449: q <= 32'b10111111010111000110110111101000 ;
        450: q <= 32'b10111111011110010101000011101001 ;
        451: q <= 32'b10111111011010010001001111010010 ;
        452: q <= 32'b00111110010010011000001111101100 ;
        453: q <= 32'b10111110100010000100010000110100 ;
        454: q <= 32'b00111110100001100010000000011111 ;
        455: q <= 32'b10111110100001001110111011100111 ;
        456: q <= 32'b10111110101010110011001100011101 ;
        457: q <= 32'b10111110010001100010100111100100 ;
        458: q <= 32'b00111110011001111011000000010111 ;
        459: q <= 32'b10111101000011100101010101110110 ;
        460: q <= 32'b00111110100110000111111110111001 ;
        461: q <= 32'b10111110100011001100110001110000 ;
        462: q <= 32'b00111101111100001010111010000010 ;
        463: q <= 32'b00111110100010100001000011101110 ;
        464: q <= 32'b10111110010000101000011000100001 ;
        465: q <= 32'b10111111001111100000111111111000 ;
        466: q <= 32'b00111110110101010100001010110110 ;
        467: q <= 32'b10111101001111110111000101111100 ;
        468: q <= 32'b00111110111101111101000001100010 ;
        469: q <= 32'b00111101100101000101010011101011 ;
        470: q <= 32'b00111110000101011110110111111101 ;
        471: q <= 32'b00111110000000100010111110001001 ;
        472: q <= 32'b00111111001010110000011011000111 ;
        473: q <= 32'b00111101010000111010110001011111 ;
        474: q <= 32'b10111110000101011101010010001000 ;
        475: q <= 32'b00111110101010111110100001100100 ;
        476: q <= 32'b00111111000001001101010011110100 ;
        477: q <= 32'b10111110100000001110001001010110 ;
        478: q <= 32'b10111101100010111000110101101001 ;
        479: q <= 32'b00111100101011001011110101010001 ;
        480: q <= 32'b10111110010000001101101110001100 ;
        481: q <= 32'b10111101100110110101110100001010 ;
        482: q <= 32'b00111111011010011001101101100110 ;
        483: q <= 32'b00111110100010110010001101100101 ;
        484: q <= 32'b00111110001011001111011111010111 ;
        485: q <= 32'b10111101000100011001111001001111 ;
        486: q <= 32'b00111101010011111010100111011100 ;
        487: q <= 32'b00111111000110011110100011101001 ;
        488: q <= 32'b10111110100011111000110101010101 ;
        489: q <= 32'b00111110100000001001001000010111 ;
        490: q <= 32'b00111110001101100111010100001000 ;
        491: q <= 32'b00111110100101111010110011111000 ;
        492: q <= 32'b10111110011011101111110100000100 ;
        493: q <= 32'b00111101110011111100101101101001 ;
        494: q <= 32'b10111110010111100110011101111000 ;
        495: q <= 32'b10111101101010001110011000010000 ;
        496: q <= 32'b00111110100001110000001011100101 ;
        497: q <= 32'b10111110101000000001101011110011 ;
        498: q <= 32'b10111110000001011001110011010110 ;
        499: q <= 32'b10111101010100111111000101011001 ;
        500: q <= 32'b00111101111101111110101100010110 ;
        501: q <= 32'b10111100111111001101000101011011 ;
        502: q <= 32'b00111110011110001101111101111101 ;
        503: q <= 32'b00111101000001110001000101010010 ;
        504: q <= 32'b00111110001000100000101010011101 ;
        505: q <= 32'b00111101000101011001100111001100 ;
        506: q <= 32'b00111110100011111101010101101111 ;
        507: q <= 32'b10111101111101000111001100110101 ;
        508: q <= 32'b00000000000000000000000000000000 ;
        509: q <= 32'b00000000000000000000000000000000 ;
        510: q <= 32'b00000000000000000000000000000000 ;
        511: q <= 32'b00000000000000000000000000000000 ;
        512: q <= 32'b00111111001000001100100000110101 ;
        513: q <= 32'b00111101100110100011101001110110 ;
        514: q <= 32'b10111101111000001101101010110110 ;
        515: q <= 32'b10111101100100110100011010000011 ;
        516: q <= 32'b10111101001100000001000101100000 ;
        517: q <= 32'b10111110000001111101010000011001 ;
        518: q <= 32'b10111101011100010000000111111011 ;
        519: q <= 32'b10111110100110110010000011001010 ;
        520: q <= 32'b00111111000110100001001010011110 ;
        521: q <= 32'b10111110100001001001111110100000 ;
        522: q <= 32'b00111101010111100001110111000001 ;
        523: q <= 32'b10111110011000001010001011001000 ;
        524: q <= 32'b10111110110010011101011010001010 ;
        525: q <= 32'b10111101101001010101001100000100 ;
        526: q <= 32'b00111110100101011101011001011011 ;
        527: q <= 32'b00111110001101010101000010101100 ;
        528: q <= 32'b10111111001001000000110010001100 ;
        529: q <= 32'b00111101100101101011001111100101 ;
        530: q <= 32'b00111110110011100110100011011101 ;
        531: q <= 32'b00111101110110100110010010101001 ;
        532: q <= 32'b10111110101100010101111010111011 ;
        533: q <= 32'b00111101110101010110010000101011 ;
        534: q <= 32'b00111101100101101100011010110111 ;
        535: q <= 32'b00111110010001111011110010000001 ;
        536: q <= 32'b10111110100110011110010011001000 ;
        537: q <= 32'b00111101110011001110010010000011 ;
        538: q <= 32'b00111111000000011010100010010000 ;
        539: q <= 32'b00111110100110101001101010101000 ;
        540: q <= 32'b10111101111110000011000010000101 ;
        541: q <= 32'b10111110101010100111000111011100 ;
        542: q <= 32'b00111101100110001101101010111011 ;
        543: q <= 32'b10111110101000001111010110101011 ;
        544: q <= 32'b10111110101111111011111000101110 ;
        545: q <= 32'b10111110001010011000110001111100 ;
        546: q <= 32'b10111110010001101010110000001010 ;
        547: q <= 32'b10111111010010011010101010011110 ;
        548: q <= 32'b00111110010000111000001110001010 ;
        549: q <= 32'b00111101011011001100011011101101 ;
        550: q <= 32'b00111101110001011111111110111101 ;
        551: q <= 32'b10111110101000010000001001001011 ;
        552: q <= 32'b10111100100110100001111100110110 ;
        553: q <= 32'b10111111001101010000110011110100 ;
        554: q <= 32'b00111101111011000010001111111111 ;
        555: q <= 32'b00111110001111110011110010011111 ;
        556: q <= 32'b10111110100111001010111010000101 ;
        557: q <= 32'b00111101010111111100011101100001 ;
        558: q <= 32'b10111110001100101000000110100111 ;
        559: q <= 32'b10111111010101100001111011110111 ;
        560: q <= 32'b00111101101111011101001011001110 ;
        561: q <= 32'b10111110010111100111111000001001 ;
        562: q <= 32'b10111110101010001101110011110011 ;
        563: q <= 32'b10111110001111100110111110101111 ;
        564: q <= 32'b10111101001110010000101111110111 ;
        565: q <= 32'b10111101011100100110011101100000 ;
        566: q <= 32'b10111111011010001110000011010011 ;
        567: q <= 32'b10111100101111100011110011010010 ;
        568: q <= 32'b00111110001100101110111111001110 ;
        569: q <= 32'b10111101100100110001101110111010 ;
        570: q <= 32'b00111110010110101011101111011100 ;
        571: q <= 32'b10111110100111000101011100000100 ;
        572: q <= 32'b00000000000000000000000000000000 ;
        573: q <= 32'b00000000000000000000000000000000 ;
        574: q <= 32'b00000000000000000000000000000000 ;
        575: q <= 32'b00000000000000000000000000000000 ;
        576: q <= 32'b10111100011100111101011000000100 ;
        577: q <= 32'b00111101111010001100110001101001 ;
        578: q <= 32'b10111101100010101101100011001111 ;
        579: q <= 32'b10111100100001110001001010100101 ;
        580: q <= 32'b00111101001010111000100100000101 ;
        581: q <= 32'b10111110001001000011110111110001 ;
        582: q <= 32'b10111100101100101011110101111010 ;
        583: q <= 32'b10111101101101011010010110111011 ;
        584: q <= 32'b00111110101100101001110010011110 ;
        585: q <= 32'b10111110001110000001011111110010 ;
        586: q <= 32'b00111110000011111100000100110100 ;
        587: q <= 32'b00111110000100110011000011011110 ;
        588: q <= 32'b10111110101001110111111011011100 ;
        589: q <= 32'b10111110010011000001011110110010 ;
        590: q <= 32'b00111101001000111111001000011001 ;
        591: q <= 32'b00111110010110000111010011110110 ;
        592: q <= 32'b00111110010100101101000001011101 ;
        593: q <= 32'b10111110111111110101010101100101 ;
        594: q <= 32'b10111110101010100001010011001001 ;
        595: q <= 32'b00111110000111101001010110111000 ;
        596: q <= 32'b00111110101001000010001100100110 ;
        597: q <= 32'b00111101101110001111110001000100 ;
        598: q <= 32'b10111101011100100111110111000001 ;
        599: q <= 32'b00111101100111100001011100101010 ;
        600: q <= 32'b00111110101110010110011011011110 ;
        601: q <= 32'b10111110101110110110101100111111 ;
        602: q <= 32'b00111110100011010101100100100010 ;
        603: q <= 32'b00111110100000110011000010111111 ;
        604: q <= 32'b10111110000011011111001010011111 ;
        605: q <= 32'b10111110010000110101000100010101 ;
        606: q <= 32'b00111101110011011001001001101011 ;
        607: q <= 32'b10111101110001011000110000111100 ;
        608: q <= 32'b00111110111000000101110101100111 ;
        609: q <= 32'b00111011111001101101111001010110 ;
        610: q <= 32'b10111110011100110100101001000100 ;
        611: q <= 32'b00111100011001111010010010100011 ;
        612: q <= 32'b00111110000000000010010111010011 ;
        613: q <= 32'b10111110010010011101110100000111 ;
        614: q <= 32'b10111111000111000111100010001010 ;
        615: q <= 32'b10111110001101011000001110011000 ;
        616: q <= 32'b10111110001100110000011010100000 ;
        617: q <= 32'b10111110010011111100011000101011 ;
        618: q <= 32'b00111100101001101101010110101000 ;
        619: q <= 32'b00111101111110101101011011101001 ;
        620: q <= 32'b10111110000010111110001100101111 ;
        621: q <= 32'b10111110000111111110100100011100 ;
        622: q <= 32'b10111111010010000101000111011010 ;
        623: q <= 32'b10111111001001101111110101101100 ;
        624: q <= 32'b00111110000110110111101010100000 ;
        625: q <= 32'b10111101110100100111001110011010 ;
        626: q <= 32'b10111110001011000100010001000000 ;
        627: q <= 32'b00111111000010001011001001101011 ;
        628: q <= 32'b00111111010010011011100011111000 ;
        629: q <= 32'b10111101010011100001100100111000 ;
        630: q <= 32'b00111110100000101011110100110100 ;
        631: q <= 32'b00111100111000000110011110110010 ;
        632: q <= 32'b00111110011010111101001000001001 ;
        633: q <= 32'b00111101111101100011111000011011 ;
        634: q <= 32'b00111101101101111000011010101011 ;
        635: q <= 32'b10111110010000110110100101101000 ;
        636: q <= 32'b00000000000000000000000000000000 ;
        637: q <= 32'b00000000000000000000000000000000 ;
        638: q <= 32'b00000000000000000000000000000000 ;
        639: q <= 32'b00000000000000000000000000000000 ;
        640: q <= 32'b10111101100001111010010100000001 ;
        641: q <= 32'b10111111010010010101100000111101 ;
        642: q <= 32'b00111101000101101111000110111001 ;
        643: q <= 32'b10111101101111111110011001010001 ;
        644: q <= 32'b00111101111110110110001100000101 ;
        645: q <= 32'b10111110100101101101101101110010 ;
        646: q <= 32'b10111110010010101000001011011000 ;
        647: q <= 32'b10111110100010000111111001001011 ;
        648: q <= 32'b10111110001010000011010111101001 ;
        649: q <= 32'b10111110010111000001010001101100 ;
        650: q <= 32'b00111101100010000100001001111000 ;
        651: q <= 32'b10111110000100111010001010110100 ;
        652: q <= 32'b00111110110100011110101111010111 ;
        653: q <= 32'b10111110001101110111111101010111 ;
        654: q <= 32'b00111110101100011101110010011011 ;
        655: q <= 32'b00111110010100111010000101010010 ;
        656: q <= 32'b00111101000001110011010111011110 ;
        657: q <= 32'b00111101011000001111111001100001 ;
        658: q <= 32'b10111111000110111110111110011111 ;
        659: q <= 32'b00111111000001001011111110011010 ;
        660: q <= 32'b00111111000011011011101100011001 ;
        661: q <= 32'b00111110101110010011001010000010 ;
        662: q <= 32'b10111110001011010001100010110010 ;
        663: q <= 32'b00111110101101100011100100001100 ;
        664: q <= 32'b00111111001001010110000000000100 ;
        665: q <= 32'b00111101110100010101101111001110 ;
        666: q <= 32'b00111111001100111000100100011001 ;
        667: q <= 32'b00111110100101100010100000111011 ;
        668: q <= 32'b00111111000110110011110010011011 ;
        669: q <= 32'b10111110100010101101010100110101 ;
        670: q <= 32'b10111101111001000001101010111100 ;
        671: q <= 32'b00111100000100111001100000010011 ;
        672: q <= 32'b00111111000111110110110001101010 ;
        673: q <= 32'b00111101001011110001101000101111 ;
        674: q <= 32'b10111110101011001110111010100111 ;
        675: q <= 32'b10111111010011010000011010011110 ;
        676: q <= 32'b00111110011010010011001110100100 ;
        677: q <= 32'b10111010100111001110000101100001 ;
        678: q <= 32'b10111110010001001010100010011100 ;
        679: q <= 32'b10111111000110110101001110010101 ;
        680: q <= 32'b10111110010110111110000010110000 ;
        681: q <= 32'b00111110111001101010001011001100 ;
        682: q <= 32'b00111101101111101000000011101001 ;
        683: q <= 32'b10111111000100001010110100000111 ;
        684: q <= 32'b10111101111010000110000010010010 ;
        685: q <= 32'b10111101110010100111010010001111 ;
        686: q <= 32'b10111101001010110011001100010110 ;
        687: q <= 32'b10111101000000101101000001010110 ;
        688: q <= 32'b10111110000011011011111001011000 ;
        689: q <= 32'b10111110100101110100101011101011 ;
        690: q <= 32'b10111110100000011100110100100101 ;
        691: q <= 32'b10111110001111000000101000001100 ;
        692: q <= 32'b10111101000101101000000011110110 ;
        693: q <= 32'b10111101101000100011110100011011 ;
        694: q <= 32'b10111111010010000010110101100010 ;
        695: q <= 32'b10111100100101100110001110000101 ;
        696: q <= 32'b00111110011100110101101011100100 ;
        697: q <= 32'b00111101111110101111100110110000 ;
        698: q <= 32'b00111110100011011000001101000010 ;
        699: q <= 32'b10111110101110101110011100110100 ;
        700: q <= 32'b00000000000000000000000000000000 ;
        701: q <= 32'b00000000000000000000000000000000 ;
        702: q <= 32'b00000000000000000000000000000000 ;
        703: q <= 32'b00000000000000000000000000000000 ;
        704: q <= 32'b10111101111011100110010000000000 ;
        705: q <= 32'b00111110111010111110101001101011 ;
        706: q <= 32'b10111111011001001001101011101100 ;
        707: q <= 32'b00111101101001001111110111111011 ;
        708: q <= 32'b00111110000010011001001101101000 ;
        709: q <= 32'b10111110010100001001100000010100 ;
        710: q <= 32'b10111110010111100011000111111110 ;
        711: q <= 32'b10111110100111010100101100100001 ;
        712: q <= 32'b00111111011100110011001111111000 ;
        713: q <= 32'b10111110100110101110111111000101 ;
        714: q <= 32'b00111100111100101100011001100011 ;
        715: q <= 32'b10111110000010100101101000100110 ;
        716: q <= 32'b10111111000010110001001001111000 ;
        717: q <= 32'b10111101111110000110101110010011 ;
        718: q <= 32'b00111101110110111001011011010001 ;
        719: q <= 32'b00111110011010010001111100100000 ;
        720: q <= 32'b00111110000110110010000101101000 ;
        721: q <= 32'b00111110101001000111011000110011 ;
        722: q <= 32'b10111110111010011101010110000111 ;
        723: q <= 32'b10111100111000001001000001101010 ;
        724: q <= 32'b00111110100010101000010011000100 ;
        725: q <= 32'b00111110000000011111111100111000 ;
        726: q <= 32'b10111101110010101101111100111001 ;
        727: q <= 32'b10111110001001010000011000110101 ;
        728: q <= 32'b00111110111000011011111010101111 ;
        729: q <= 32'b10111101001110010111111101001010 ;
        730: q <= 32'b10111110101100010001001000000000 ;
        731: q <= 32'b00111110011101101110110001001110 ;
        732: q <= 32'b00111111000000010010111001110111 ;
        733: q <= 32'b10111110101010110001000011011001 ;
        734: q <= 32'b00111111100010011111111011011011 ;
        735: q <= 32'b00111101110011011100110011101001 ;
        736: q <= 32'b10111101110110100011001111001111 ;
        737: q <= 32'b00111101110101011001011111110100 ;
        738: q <= 32'b10111110101011111101100101101010 ;
        739: q <= 32'b00111011011001100000001110010000 ;
        740: q <= 32'b00111110011101000110010110010011 ;
        741: q <= 32'b00111110010110010011100100100010 ;
        742: q <= 32'b10111101000010100110011110010100 ;
        743: q <= 32'b00111110110110100110111010000000 ;
        744: q <= 32'b10111101100100100001110000110100 ;
        745: q <= 32'b00111110100011100100011101000000 ;
        746: q <= 32'b00111101101011010101100000011101 ;
        747: q <= 32'b00111110001010011000001110100110 ;
        748: q <= 32'b10111110101000110011111001100100 ;
        749: q <= 32'b10111100111000011110111111000011 ;
        750: q <= 32'b10111011110001010011101001000001 ;
        751: q <= 32'b00111011000101110000010000110000 ;
        752: q <= 32'b00111110011010010000111011111011 ;
        753: q <= 32'b10111110101000011110000111110010 ;
        754: q <= 32'b10111110100011111001011111100100 ;
        755: q <= 32'b10111110000010100100111000010011 ;
        756: q <= 32'b10111011101010000000011111000000 ;
        757: q <= 32'b00111101110100011000101101110100 ;
        758: q <= 32'b10111111010100011001101011011010 ;
        759: q <= 32'b00111110000000011011000111001010 ;
        760: q <= 32'b00111110100100100011001010111011 ;
        761: q <= 32'b10111101000100110010111001001010 ;
        762: q <= 32'b00111101011110100110111110101110 ;
        763: q <= 32'b10111110011010000110000011110101 ;
        764: q <= 32'b00000000000000000000000000000000 ;
        765: q <= 32'b00000000000000000000000000000000 ;
        766: q <= 32'b00000000000000000000000000000000 ;
        767: q <= 32'b00000000000000000000000000000000 ;
        768: q <= 32'b10111110001011110010010001111011 ;
        769: q <= 32'b00111110000101000100111110110100 ;
        770: q <= 32'b00111110000110001110101010000100 ;
        771: q <= 32'b10111110100011001000100101011011 ;
        772: q <= 32'b10111101000010100000111010110110 ;
        773: q <= 32'b10111110101110001110110110011110 ;
        774: q <= 32'b00111110010010110000101111011000 ;
        775: q <= 32'b10111110000010101100111011111011 ;
        776: q <= 32'b10111101110110001010010100011011 ;
        777: q <= 32'b10111110011001111100000110101110 ;
        778: q <= 32'b00111110010001101111010011100100 ;
        779: q <= 32'b10111110000011110010001011000001 ;
        780: q <= 32'b10111110100011101000111101101101 ;
        781: q <= 32'b10111110100100011000110000101111 ;
        782: q <= 32'b00111101110011111011001001010011 ;
        783: q <= 32'b00111110010100101010101001010100 ;
        784: q <= 32'b10111111001000011110101000001000 ;
        785: q <= 32'b00111101001101010100000101010111 ;
        786: q <= 32'b10111110111000010111111001111111 ;
        787: q <= 32'b00111110010010100000000101000111 ;
        788: q <= 32'b10111110101011100000010000110111 ;
        789: q <= 32'b00111110000110001000010010101111 ;
        790: q <= 32'b00111111011100100101100100001110 ;
        791: q <= 32'b00111111011001000010111011001100 ;
        792: q <= 32'b00111110101110110000100111111011 ;
        793: q <= 32'b10111110001010101100000110010111 ;
        794: q <= 32'b10111110110110001011011100101011 ;
        795: q <= 32'b00111110000001110000010100010111 ;
        796: q <= 32'b00111111001000111010000001111000 ;
        797: q <= 32'b10111110101000110111010101110010 ;
        798: q <= 32'b00111011111100001010111000101111 ;
        799: q <= 32'b00111101101001010010101100110010 ;
        800: q <= 32'b00111110000101110111001010000000 ;
        801: q <= 32'b10111111100000110110111001001011 ;
        802: q <= 32'b10111110110100101111101010010000 ;
        803: q <= 32'b00111101110001111101111010101110 ;
        804: q <= 32'b00111110010111001110110000010101 ;
        805: q <= 32'b10111101001011110000111000101100 ;
        806: q <= 32'b10111101100110001110110000101110 ;
        807: q <= 32'b00111110100111110101101001011100 ;
        808: q <= 32'b10111110100111001010011101110111 ;
        809: q <= 32'b00111110011011010011001011110100 ;
        810: q <= 32'b00111100110001011100000111010001 ;
        811: q <= 32'b00111110001010011011001110100100 ;
        812: q <= 32'b10111110001110100101101001010010 ;
        813: q <= 32'b00111101110010001101111011111011 ;
        814: q <= 32'b10111110100110010011111011101110 ;
        815: q <= 32'b10111101011100111110001101101111 ;
        816: q <= 32'b10111111001110110000000111111111 ;
        817: q <= 32'b10111110011111010110001010000001 ;
        818: q <= 32'b10111110101000111001101000110101 ;
        819: q <= 32'b10111101110101110011010100100101 ;
        820: q <= 32'b00111110100011011111001011000001 ;
        821: q <= 32'b00111101000010111100101111011011 ;
        822: q <= 32'b00111110010001110100100011111011 ;
        823: q <= 32'b10111101101000110101100001100011 ;
        824: q <= 32'b00111110100101110000001011100001 ;
        825: q <= 32'b10111101100001100001010011101000 ;
        826: q <= 32'b00111110010001101100001001110000 ;
        827: q <= 32'b10111110010000110111001000001100 ;
        828: q <= 32'b00000000000000000000000000000000 ;
        829: q <= 32'b00000000000000000000000000000000 ;
        830: q <= 32'b00000000000000000000000000000000 ;
        831: q <= 32'b00000000000000000000000000000000 ;
        832: q <= 32'b00111101100111110111001011111010 ;
        833: q <= 32'b00111110001000100010010001101111 ;
        834: q <= 32'b00111100100110010001010011111111 ;
        835: q <= 32'b10111101101101001100011001011101 ;
        836: q <= 32'b00111110000010111010010101100101 ;
        837: q <= 32'b10111101101011110010010010011111 ;
        838: q <= 32'b10111111000111101011100111000001 ;
        839: q <= 32'b10111110100110100111100111011000 ;
        840: q <= 32'b00111101101100010010001101111110 ;
        841: q <= 32'b10111110000001001000100010110010 ;
        842: q <= 32'b00111110100000010110101000110010 ;
        843: q <= 32'b10111111001100111100110000000010 ;
        844: q <= 32'b00111110101111111001011110101110 ;
        845: q <= 32'b10111101101101000011101111001001 ;
        846: q <= 32'b00111110001011110100001000001110 ;
        847: q <= 32'b00111110100010110000001010000010 ;
        848: q <= 32'b00111110100000101100101110010011 ;
        849: q <= 32'b10111110111000100111101110110010 ;
        850: q <= 32'b10111110100001111101101000111010 ;
        851: q <= 32'b00111110011001100101011101101111 ;
        852: q <= 32'b10111110101101000010111101101100 ;
        853: q <= 32'b00111110000101001010111001001110 ;
        854: q <= 32'b00111110101110000100100111111111 ;
        855: q <= 32'b00111110000110100010010011100001 ;
        856: q <= 32'b00111110111010101001001011010110 ;
        857: q <= 32'b00111110001100111100011100100100 ;
        858: q <= 32'b00111110100110011100101010001100 ;
        859: q <= 32'b00111110001100011010001110110111 ;
        860: q <= 32'b10111100111111010011001001000100 ;
        861: q <= 32'b10111101111100000010011000000111 ;
        862: q <= 32'b00111110001010000100011010101001 ;
        863: q <= 32'b10111101010111001110111001100011 ;
        864: q <= 32'b10111110010011010010100100001101 ;
        865: q <= 32'b10111101011001011100101000001011 ;
        866: q <= 32'b10111110100110111000101011111010 ;
        867: q <= 32'b10111101101110010101000000111011 ;
        868: q <= 32'b10111100001000011011100110011100 ;
        869: q <= 32'b10111110110010111100010110000011 ;
        870: q <= 32'b00111101101110001000101000011010 ;
        871: q <= 32'b00111111000101011000010000110001 ;
        872: q <= 32'b10111110011001001011100111000111 ;
        873: q <= 32'b10111110110010111100101010000110 ;
        874: q <= 32'b00111111001110110100111001101101 ;
        875: q <= 32'b10111110100010000011000010101010 ;
        876: q <= 32'b10111110101000100011101100011110 ;
        877: q <= 32'b10111101101110110010011100100010 ;
        878: q <= 32'b10111110011001101000010000010101 ;
        879: q <= 32'b10111101110101111100011011011111 ;
        880: q <= 32'b00111110100010001100000010001101 ;
        881: q <= 32'b10111110101011000100001101010101 ;
        882: q <= 32'b10111110010001100000000111001110 ;
        883: q <= 32'b10111110100111110101011001011101 ;
        884: q <= 32'b00111101100100100111101101001110 ;
        885: q <= 32'b00111111000010110110100110111000 ;
        886: q <= 32'b00111101010011000100001000000110 ;
        887: q <= 32'b00111111001001001010110011010001 ;
        888: q <= 32'b00111110100011100101011110001100 ;
        889: q <= 32'b10111111000010111001011111100100 ;
        890: q <= 32'b00111110001110000010100110011010 ;
        891: q <= 32'b10111110011111110000101111100001 ;
        892: q <= 32'b00000000000000000000000000000000 ;
        893: q <= 32'b00000000000000000000000000000000 ;
        894: q <= 32'b00000000000000000000000000000000 ;
        895: q <= 32'b00000000000000000000000000000000 ;
        896: q <= 32'b00111111000110000101111110101110 ;
        897: q <= 32'b00111110010110000000000010011001 ;
        898: q <= 32'b10111101100101101011001010111101 ;
        899: q <= 32'b10111101001111100011111001010001 ;
        900: q <= 32'b00111101110111110000111110110010 ;
        901: q <= 32'b10111110101011111101011110111001 ;
        902: q <= 32'b10111110000101101110001001101110 ;
        903: q <= 32'b10111110101110010111101100101000 ;
        904: q <= 32'b00111111011001100000100000101010 ;
        905: q <= 32'b10111110100100001111000010110111 ;
        906: q <= 32'b00111110101101010100001101000100 ;
        907: q <= 32'b10111110001001110110010101001011 ;
        908: q <= 32'b00111111000101100000101001000101 ;
        909: q <= 32'b10111110100110010101000110000001 ;
        910: q <= 32'b10111111010100010010111010001000 ;
        911: q <= 32'b00111110100001000010111100100101 ;
        912: q <= 32'b00111110001001111100000110001010 ;
        913: q <= 32'b00111100111001011110011001110001 ;
        914: q <= 32'b00111101111100110100001001100101 ;
        915: q <= 32'b00111100010110101100100100101001 ;
        916: q <= 32'b10111110110101100100111100000000 ;
        917: q <= 32'b00111110100010010100110000000100 ;
        918: q <= 32'b00111100100110011111010100010010 ;
        919: q <= 32'b00111101101101100100011000110000 ;
        920: q <= 32'b10111110010011101000000100000100 ;
        921: q <= 32'b00111110011111111000001100011111 ;
        922: q <= 32'b10111110100111000111101001010101 ;
        923: q <= 32'b00111110100111111101101000011100 ;
        924: q <= 32'b10111101000110100110010110101000 ;
        925: q <= 32'b10111111001001001000101011101010 ;
        926: q <= 32'b00111110001000100111111010100010 ;
        927: q <= 32'b10111111010001001101110001110110 ;
        928: q <= 32'b00111111011100010001110010101000 ;
        929: q <= 32'b10111101101010010001011100000001 ;
        930: q <= 32'b10111110010000101011000111000011 ;
        931: q <= 32'b00111110100000100111100100011001 ;
        932: q <= 32'b00111110100101111101011111100110 ;
        933: q <= 32'b00111100100010101010011111010110 ;
        934: q <= 32'b00111100100110001000111011010001 ;
        935: q <= 32'b10111110111101001111101100000001 ;
        936: q <= 32'b10111010111010000100001111100110 ;
        937: q <= 32'b00111110101101010101001001101010 ;
        938: q <= 32'b10111101010100111011011110001101 ;
        939: q <= 32'b00111111001010001001101111000111 ;
        940: q <= 32'b10111110101001110111111101000011 ;
        941: q <= 32'b10111100011000110110110111011110 ;
        942: q <= 32'b10111110000111000101100111101101 ;
        943: q <= 32'b00111101001000010100100100011000 ;
        944: q <= 32'b00111110101101000010110010011110 ;
        945: q <= 32'b10111110110010000010011001001101 ;
        946: q <= 32'b10111110101011000111001010000101 ;
        947: q <= 32'b10111110011011100000010110000011 ;
        948: q <= 32'b00111110010110011110010101100101 ;
        949: q <= 32'b00111100010011111111001001000010 ;
        950: q <= 32'b00111110110011111111100110111011 ;
        951: q <= 32'b00111110010000010100101000101110 ;
        952: q <= 32'b00111110101101110010100011110111 ;
        953: q <= 32'b10111101011001100000100101010111 ;
        954: q <= 32'b00111110010011001011001100001001 ;
        955: q <= 32'b10111110110101000011110110101011 ;
        956: q <= 32'b00000000000000000000000000000000 ;
        957: q <= 32'b00000000000000000000000000000000 ;
        958: q <= 32'b00000000000000000000000000000000 ;
        959: q <= 32'b00000000000000000000000000000000 ;
        960: q <= 32'b10111110000011101110001000101011 ;
        961: q <= 32'b00111110000000110001010110100010 ;
        962: q <= 32'b00111101011010111000001000110000 ;
        963: q <= 32'b10111111011101000111010111111000 ;
        964: q <= 32'b00111110001001000111000011011011 ;
        965: q <= 32'b10111110100010000011101010010000 ;
        966: q <= 32'b10111111011000111010011010100011 ;
        967: q <= 32'b10111110011001010010111111011011 ;
        968: q <= 32'b10111101100111100111000101100100 ;
        969: q <= 32'b10111110101001101010000001000111 ;
        970: q <= 32'b10111111001000110001001000011011 ;
        971: q <= 32'b00111110010011011100101001000100 ;
        972: q <= 32'b00111110110001100011100110000001 ;
        973: q <= 32'b10111110100101101101111010000101 ;
        974: q <= 32'b00111110011000000011110101100100 ;
        975: q <= 32'b00111110100110110010100100010101 ;
        976: q <= 32'b00111110110000000011100111100100 ;
        977: q <= 32'b10111111010000000000010111011101 ;
        978: q <= 32'b00111111000101101110011101001110 ;
        979: q <= 32'b00111110000001001110111111110010 ;
        980: q <= 32'b10111110110110100011111100000101 ;
        981: q <= 32'b00111101111110010101110001110011 ;
        982: q <= 32'b10111110001100110111001111001101 ;
        983: q <= 32'b00111110100100000111011110111010 ;
        984: q <= 32'b10111110111000001001001111111111 ;
        985: q <= 32'b00111101100011011101000001100101 ;
        986: q <= 32'b10111111000101101101011101101100 ;
        987: q <= 32'b00111110101011101101101110111101 ;
        988: q <= 32'b10111110000011100111010110100000 ;
        989: q <= 32'b10111110100011010001111110010110 ;
        990: q <= 32'b00111110100010000101011101000000 ;
        991: q <= 32'b00111101010001010001110110010101 ;
        992: q <= 32'b00111111000011110000010111110000 ;
        993: q <= 32'b10111101001101111110000010111100 ;
        994: q <= 32'b00111110111001101100101101111000 ;
        995: q <= 32'b10111110010000101110111011001001 ;
        996: q <= 32'b10111100011011110110101110011010 ;
        997: q <= 32'b10111101010101110001000110100011 ;
        998: q <= 32'b00111110000011011100010000011110 ;
        999: q <= 32'b10111110100100110110111010001001 ;
        1000: q <= 32'b00111100011011000111011110110000 ;
        1001: q <= 32'b10111111000100111011000000110000 ;
        1002: q <= 32'b00111100011011010000111011001011 ;
        1003: q <= 32'b10111110100011110011000000111111 ;
        1004: q <= 32'b10111110010010110100010100000010 ;
        1005: q <= 32'b00111110100100010010000110000011 ;
        1006: q <= 32'b10111101110110000010101011111100 ;
        1007: q <= 32'b10111110010010000110011111011111 ;
        1008: q <= 32'b10111101000111100001101000011010 ;
        1009: q <= 32'b10111110101100010011110111001101 ;
        1010: q <= 32'b10111110000010110000010001110100 ;
        1011: q <= 32'b00111111000100100011110011011101 ;
        1012: q <= 32'b00111100101001001001000111000100 ;
        1013: q <= 32'b10111101100110111100001000100001 ;
        1014: q <= 32'b00111101001100101110011010000000 ;
        1015: q <= 32'b00111101100110010110001000000100 ;
        1016: q <= 32'b00111110011111011011011111001111 ;
        1017: q <= 32'b00111110001001011100100010000111 ;
        1018: q <= 32'b00111110100011110000000000111011 ;
        1019: q <= 32'b10111110100010110010101010011001 ;
        1020: q <= 32'b00000000000000000000000000000000 ;
        1021: q <= 32'b00000000000000000000000000000000 ;
        1022: q <= 32'b00000000000000000000000000000000 ;
        1023: q <= 32'b00000000000000000000000000000000 ;
        1024: q <= 32'b10111110001000011100010011110001 ;
        1025: q <= 32'b10111111010011100111111111001011 ;
        1026: q <= 32'b10111110000011001010001110010100 ;
        1027: q <= 32'b00111101110010101110111110001000 ;
        1028: q <= 32'b00111110010111101101011011010000 ;
        1029: q <= 32'b10111101111110110000010001001011 ;
        1030: q <= 32'b10111111010010100110001011111010 ;
        1031: q <= 32'b10111110100111011011111011001010 ;
        1032: q <= 32'b00111011100101011100101101101111 ;
        1033: q <= 32'b10111101011100001001011110110001 ;
        1034: q <= 32'b00111110110110011101100001100111 ;
        1035: q <= 32'b10111100101001111100101110001011 ;
        1036: q <= 32'b10111110100010011010011000010100 ;
        1037: q <= 32'b10111110010110101101111000010010 ;
        1038: q <= 32'b10111110101110000101111011011110 ;
        1039: q <= 32'b00111110001111111000011111110101 ;
        1040: q <= 32'b10111111000110011000000001001010 ;
        1041: q <= 32'b00111110010011100011001010011010 ;
        1042: q <= 32'b00111111000011011110100000010010 ;
        1043: q <= 32'b00111111000010110001001100100100 ;
        1044: q <= 32'b00111111010001100011100000011111 ;
        1045: q <= 32'b00111110001100000110110000001110 ;
        1046: q <= 32'b00111110000100101001100101000000 ;
        1047: q <= 32'b00111110100000101110001110111101 ;
        1048: q <= 32'b10111110001101100000000101101001 ;
        1049: q <= 32'b10111100000110010010010101001110 ;
        1050: q <= 32'b10111110100000010110110100011011 ;
        1051: q <= 32'b00111110100111111010111011110001 ;
        1052: q <= 32'b00111100100101011001111011111011 ;
        1053: q <= 32'b10111110000011111011110101010110 ;
        1054: q <= 32'b00111101101010101101101110011000 ;
        1055: q <= 32'b10111101100011001110101001110111 ;
        1056: q <= 32'b10111101101010001101000010110011 ;
        1057: q <= 32'b00111110010000101101101001100111 ;
        1058: q <= 32'b10111111000011101111111101110000 ;
        1059: q <= 32'b00111101100100111000000110000010 ;
        1060: q <= 32'b00111101101010110100011000000011 ;
        1061: q <= 32'b00111111000111011111111011101011 ;
        1062: q <= 32'b10111101111101100111001001111010 ;
        1063: q <= 32'b00111110101010010111000101111111 ;
        1064: q <= 32'b00111100010000100001101010011001 ;
        1065: q <= 32'b10111110111011010100100110100011 ;
        1066: q <= 32'b10111101001111111111110111010000 ;
        1067: q <= 32'b00111110100101101001011001101101 ;
        1068: q <= 32'b10111110001010011110011110011000 ;
        1069: q <= 32'b10111111010000001001101010000000 ;
        1070: q <= 32'b10111110100000000110000010010000 ;
        1071: q <= 32'b10111101101000101010001000111101 ;
        1072: q <= 32'b00111110000001101011000010000101 ;
        1073: q <= 32'b10111110000000100010010010111100 ;
        1074: q <= 32'b10111101101010000110001101111011 ;
        1075: q <= 32'b10111101010010000100011011010110 ;
        1076: q <= 32'b00111110011110010001001001101101 ;
        1077: q <= 32'b00111111011011011011010010010000 ;
        1078: q <= 32'b00111100000110111101110101100111 ;
        1079: q <= 32'b10111110000000100100010110110101 ;
        1080: q <= 32'b00111110011101101101011110011011 ;
        1081: q <= 32'b00111101111110001010100011101110 ;
        1082: q <= 32'b00111101110000010101001101001010 ;
        1083: q <= 32'b10111110011101111101100110001011 ;
        1084: q <= 32'b00000000000000000000000000000000 ;
        1085: q <= 32'b00000000000000000000000000000000 ;
        1086: q <= 32'b00000000000000000000000000000000 ;
        1087: q <= 32'b00000000000000000000000000000000 ;
        1088: q <= 32'b00111110110111101110100000101100 ;
        1089: q <= 32'b00111100011101010011111111000111 ;
        1090: q <= 32'b10111101100111001101010100011101 ;
        1091: q <= 32'b00111101001101011101101110101110 ;
        1092: q <= 32'b00111111100001111010110000000101 ;
        1093: q <= 32'b10111110100010001000100010000101 ;
        1094: q <= 32'b10111110111111110011101011111010 ;
        1095: q <= 32'b10111110100010010010100001100001 ;
        1096: q <= 32'b10111110101010011001011011001111 ;
        1097: q <= 32'b10111101110001101101001111100101 ;
        1098: q <= 32'b00111110110001001010011100100001 ;
        1099: q <= 32'b00111100111011000001010110010101 ;
        1100: q <= 32'b10111111000101101110110010010100 ;
        1101: q <= 32'b10111110010110001101011111110101 ;
        1102: q <= 32'b00111110010111010110011111101001 ;
        1103: q <= 32'b00111110011110001101011011110101 ;
        1104: q <= 32'b10111111001110010011010101111100 ;
        1105: q <= 32'b00111101011101000010011111100100 ;
        1106: q <= 32'b00111110111001101001000101111010 ;
        1107: q <= 32'b00111110000100101110101000111110 ;
        1108: q <= 32'b10111110111100011010111010001010 ;
        1109: q <= 32'b00111110001110110110011100111001 ;
        1110: q <= 32'b10111110000111000001100001001101 ;
        1111: q <= 32'b10111101010101110001000111000001 ;
        1112: q <= 32'b00111111001111000010010101010110 ;
        1113: q <= 32'b10111100111111101000010001011011 ;
        1114: q <= 32'b10111110100001110001010010011010 ;
        1115: q <= 32'b00111110011011111010101011010011 ;
        1116: q <= 32'b00111010010001011000010010100010 ;
        1117: q <= 32'b10111110011001111111111001101110 ;
        1118: q <= 32'b00111110001010100101101111110010 ;
        1119: q <= 32'b10111111001101111011111101010110 ;
        1120: q <= 32'b10111101001101011000001100111001 ;
        1121: q <= 32'b00111101110010010001001101011010 ;
        1122: q <= 32'b00111111000000101011001111000111 ;
        1123: q <= 32'b00111101100010100011000101100010 ;
        1124: q <= 32'b00111101100011100110110110100010 ;
        1125: q <= 32'b00111110010100001111101001111010 ;
        1126: q <= 32'b10111110110110000001101111011011 ;
        1127: q <= 32'b10111110101010001110000001101000 ;
        1128: q <= 32'b10111110000011001101101010000100 ;
        1129: q <= 32'b00111110011101010100101100010010 ;
        1130: q <= 32'b00111110010011000110110001101001 ;
        1131: q <= 32'b10111111000111001000111101001100 ;
        1132: q <= 32'b10111110000100010101110011101111 ;
        1133: q <= 32'b00111110100001101001111000000010 ;
        1134: q <= 32'b10111101111101100010110010011011 ;
        1135: q <= 32'b10111011111001000001010100110000 ;
        1136: q <= 32'b10111110010110110001111000110110 ;
        1137: q <= 32'b10111110000101100100100011010000 ;
        1138: q <= 32'b10111110100011001101110110000010 ;
        1139: q <= 32'b10111110001110101011000000001000 ;
        1140: q <= 32'b00111110010010000000010011010110 ;
        1141: q <= 32'b10111101000001011101001000010111 ;
        1142: q <= 32'b00111110101001000101100011111011 ;
        1143: q <= 32'b00111101111011000100001000101100 ;
        1144: q <= 32'b00111110010100100101111111000011 ;
        1145: q <= 32'b10111101101011001001111101110001 ;
        1146: q <= 32'b00111110010000100010011111000010 ;
        1147: q <= 32'b10111110101000010101000010110101 ;
        1148: q <= 32'b00000000000000000000000000000000 ;
        1149: q <= 32'b00000000000000000000000000000000 ;
        1150: q <= 32'b00000000000000000000000000000000 ;
        1151: q <= 32'b00000000000000000000000000000000 ;
        1152: q <= 32'b10111101101011010010101111010101 ;
        1153: q <= 32'b10111110111110000110111101110011 ;
        1154: q <= 32'b10111110010111101100001101100000 ;
        1155: q <= 32'b10111011101111100010101101010110 ;
        1156: q <= 32'b00111110000001111111011110101001 ;
        1157: q <= 32'b10111110100011101100101101011010 ;
        1158: q <= 32'b00111101101010000011111010101111 ;
        1159: q <= 32'b10111110000000011000010110011000 ;
        1160: q <= 32'b00111101010111011011011000100000 ;
        1161: q <= 32'b10111101101110100011000001000111 ;
        1162: q <= 32'b00111110010000001101000101101101 ;
        1163: q <= 32'b00111110010001000111011010111010 ;
        1164: q <= 32'b00111110101001110010111011010010 ;
        1165: q <= 32'b10111101101010000111110010101011 ;
        1166: q <= 32'b10111110001111101111101000000111 ;
        1167: q <= 32'b00111110011011100010000010101100 ;
        1168: q <= 32'b00111101011101011001011101111011 ;
        1169: q <= 32'b10111111000000100011001010101011 ;
        1170: q <= 32'b00111110101111100000001011000111 ;
        1171: q <= 32'b00111101100010101111011100001100 ;
        1172: q <= 32'b10111110111000111011011100101000 ;
        1173: q <= 32'b00111110100000010011100011100110 ;
        1174: q <= 32'b00111111000111110101100001010111 ;
        1175: q <= 32'b00111110101000011010110110001011 ;
        1176: q <= 32'b10111110101111110111000010111011 ;
        1177: q <= 32'b10111111000100011001110001001000 ;
        1178: q <= 32'b00111110101010000011100011010101 ;
        1179: q <= 32'b00111110101000001000001010100110 ;
        1180: q <= 32'b00111100101001011001010101101101 ;
        1181: q <= 32'b10111110101000100000100100110001 ;
        1182: q <= 32'b00111101110100001011001001001101 ;
        1183: q <= 32'b00111110001111001010010011101100 ;
        1184: q <= 32'b10111110001000010000101110000100 ;
        1185: q <= 32'b10111101010010100101101111101110 ;
        1186: q <= 32'b10111110011101111100100010001110 ;
        1187: q <= 32'b10111101100011110001001011101001 ;
        1188: q <= 32'b00111110001100100100001110001111 ;
        1189: q <= 32'b00111111011001111111100101010100 ;
        1190: q <= 32'b10111111001000101011110000010001 ;
        1191: q <= 32'b10111110011001000011000111010110 ;
        1192: q <= 32'b10111110000110100000010111100001 ;
        1193: q <= 32'b00111110101100110010101111011000 ;
        1194: q <= 32'b00111111001000111100001100001101 ;
        1195: q <= 32'b00111110101100110010001100100101 ;
        1196: q <= 32'b10111110000010101111101100000100 ;
        1197: q <= 32'b10111100001000100000111110111110 ;
        1198: q <= 32'b10111010100010101111010000001011 ;
        1199: q <= 32'b10111101111000110010000011111001 ;
        1200: q <= 32'b10111100000101001011010000000100 ;
        1201: q <= 32'b10111110101011011011110001001000 ;
        1202: q <= 32'b10111110011001011101101011101110 ;
        1203: q <= 32'b10111101001101001000100011010011 ;
        1204: q <= 32'b00111101111110010001101010111100 ;
        1205: q <= 32'b10111110100100010101011110110110 ;
        1206: q <= 32'b10111100110011110101111111000001 ;
        1207: q <= 32'b10111100110001000101010100000100 ;
        1208: q <= 32'b00111110000111010000101010101001 ;
        1209: q <= 32'b10111111000100101100101100111010 ;
        1210: q <= 32'b00111110001111101011101101111111 ;
        1211: q <= 32'b10111110001011000111100000110110 ;
        1212: q <= 32'b00000000000000000000000000000000 ;
        1213: q <= 32'b00000000000000000000000000000000 ;
        1214: q <= 32'b00000000000000000000000000000000 ;
        1215: q <= 32'b00000000000000000000000000000000 ;
        1216: q <= 32'b10111110001101010011001000011010 ;
        1217: q <= 32'b00111101001100010011101010101010 ;
        1218: q <= 32'b10111101100101011100101000011101 ;
        1219: q <= 32'b10111101011010011001001110111010 ;
        1220: q <= 32'b00111101001110010110100001101001 ;
        1221: q <= 32'b10111101111010011010110011101101 ;
        1222: q <= 32'b00111101101101100010011000010001 ;
        1223: q <= 32'b10111110001010111111100100000011 ;
        1224: q <= 32'b10111101110011001100000010001110 ;
        1225: q <= 32'b10111110000111101000110110110110 ;
        1226: q <= 32'b10111110101110000101110101100101 ;
        1227: q <= 32'b00111110000001111100011000000000 ;
        1228: q <= 32'b10111110011100100001111001000110 ;
        1229: q <= 32'b10111100101011000110110100001111 ;
        1230: q <= 32'b10111110110011010111110110000100 ;
        1231: q <= 32'b00111110011000100110010000100111 ;
        1232: q <= 32'b00111110010010111100010100001000 ;
        1233: q <= 32'b00111101011001101111101000011111 ;
        1234: q <= 32'b00111110100100101111100001110010 ;
        1235: q <= 32'b00111101101000101011101101111000 ;
        1236: q <= 32'b00111110101001110001001001111110 ;
        1237: q <= 32'b00111101010110001101011001111000 ;
        1238: q <= 32'b10111101100001100110001011111010 ;
        1239: q <= 32'b00111101110010100000010111101101 ;
        1240: q <= 32'b10111110011100011010001010010100 ;
        1241: q <= 32'b10111111000001101011000001011001 ;
        1242: q <= 32'b10111110100111010011100010001100 ;
        1243: q <= 32'b00111101111100101000111111011000 ;
        1244: q <= 32'b00111101100011011010010100101101 ;
        1245: q <= 32'b10111101100000111101110100101000 ;
        1246: q <= 32'b00111110001011110110011010001111 ;
        1247: q <= 32'b10111111000101001011111000001100 ;
        1248: q <= 32'b00111110101101110011001001100010 ;
        1249: q <= 32'b10111111001001001110101100111101 ;
        1250: q <= 32'b10111101111100101000101110111110 ;
        1251: q <= 32'b10111110000101010111101000011000 ;
        1252: q <= 32'b00111110000101010010001101111100 ;
        1253: q <= 32'b10111101101100011011111111100001 ;
        1254: q <= 32'b10111101101101111010000011101011 ;
        1255: q <= 32'b10111110010100100001010111011010 ;
        1256: q <= 32'b10111111001110111001000100000011 ;
        1257: q <= 32'b00111110000011111111000010000111 ;
        1258: q <= 32'b00111111000100011100100101010011 ;
        1259: q <= 32'b10111110111010011000100001110100 ;
        1260: q <= 32'b10111101101101001111100101111000 ;
        1261: q <= 32'b00111100111110011011000101100100 ;
        1262: q <= 32'b10111101011001110111100001010001 ;
        1263: q <= 32'b10111110100010001100001111101110 ;
        1264: q <= 32'b00111101111011000100100011100110 ;
        1265: q <= 32'b10111101110010011000011010010100 ;
        1266: q <= 32'b10111110000101100100000010001111 ;
        1267: q <= 32'b10111101000101101000011100010001 ;
        1268: q <= 32'b00111100010111100111011101111100 ;
        1269: q <= 32'b00111111001000101000010110011111 ;
        1270: q <= 32'b10111111000011010111001111100101 ;
        1271: q <= 32'b00111101100101001101011001001000 ;
        1272: q <= 32'b00111110011010010100100110000010 ;
        1273: q <= 32'b10111110101101101010001101001111 ;
        1274: q <= 32'b00111110010011010111100101011101 ;
        1275: q <= 32'b10111110001001110001001111100111 ;
        1276: q <= 32'b00000000000000000000000000000000 ;
        1277: q <= 32'b00000000000000000000000000000000 ;
        1278: q <= 32'b00000000000000000000000000000000 ;
        1279: q <= 32'b00000000000000000000000000000000 ;
        1280: q <= 32'b00000000000000000000000000000000 ;
        1281: q <= 32'b00000000000000000000000000000000 ;
        1282: q <= 32'b00000000000000000000000000000000 ;
        1283: q <= 32'b00000000000000000000000000000000 ;
        1284: q <= 32'b00000000000000000000000000000000 ;
        1285: q <= 32'b00000000000000000000000000000000 ;
        1286: q <= 32'b00000000000000000000000000000000 ;
        1287: q <= 32'b00000000000000000000000000000000 ;
        1288: q <= 32'b00000000000000000000000000000000 ;
        1289: q <= 32'b00000000000000000000000000000000 ;
        1290: q <= 32'b00000000000000000000000000000000 ;
        1291: q <= 32'b00000000000000000000000000000000 ;
        1292: q <= 32'b00000000000000000000000000000000 ;
        1293: q <= 32'b00000000000000000000000000000000 ;
        1294: q <= 32'b00000000000000000000000000000000 ;
        1295: q <= 32'b00000000000000000000000000000000 ;
        1296: q <= 32'b00000000000000000000000000000000 ;
        1297: q <= 32'b00000000000000000000000000000000 ;
        1298: q <= 32'b00000000000000000000000000000000 ;
        1299: q <= 32'b00000000000000000000000000000000 ;
        1300: q <= 32'b00000000000000000000000000000000 ;
        1301: q <= 32'b00000000000000000000000000000000 ;
        1302: q <= 32'b00000000000000000000000000000000 ;
        1303: q <= 32'b00000000000000000000000000000000 ;
        1304: q <= 32'b00000000000000000000000000000000 ;
        1305: q <= 32'b00000000000000000000000000000000 ;
        1306: q <= 32'b00000000000000000000000000000000 ;
        1307: q <= 32'b00000000000000000000000000000000 ;
        1308: q <= 32'b00000000000000000000000000000000 ;
        1309: q <= 32'b00000000000000000000000000000000 ;
        1310: q <= 32'b00000000000000000000000000000000 ;
        1311: q <= 32'b00000000000000000000000000000000 ;
        1312: q <= 32'b00000000000000000000000000000000 ;
        1313: q <= 32'b00000000000000000000000000000000 ;
        1314: q <= 32'b00000000000000000000000000000000 ;
        1315: q <= 32'b00000000000000000000000000000000 ;
        1316: q <= 32'b00000000000000000000000000000000 ;
        1317: q <= 32'b00000000000000000000000000000000 ;
        1318: q <= 32'b00000000000000000000000000000000 ;
        1319: q <= 32'b00000000000000000000000000000000 ;
        1320: q <= 32'b00000000000000000000000000000000 ;
        1321: q <= 32'b00000000000000000000000000000000 ;
        1322: q <= 32'b00000000000000000000000000000000 ;
        1323: q <= 32'b00000000000000000000000000000000 ;
        1324: q <= 32'b00000000000000000000000000000000 ;
        1325: q <= 32'b00000000000000000000000000000000 ;
        1326: q <= 32'b00000000000000000000000000000000 ;
        1327: q <= 32'b00000000000000000000000000000000 ;
        1328: q <= 32'b00000000000000000000000000000000 ;
        1329: q <= 32'b00000000000000000000000000000000 ;
        1330: q <= 32'b00000000000000000000000000000000 ;
        1331: q <= 32'b00000000000000000000000000000000 ;
        1332: q <= 32'b00000000000000000000000000000000 ;
        1333: q <= 32'b00000000000000000000000000000000 ;
        1334: q <= 32'b00000000000000000000000000000000 ;
        1335: q <= 32'b00000000000000000000000000000000 ;
        1336: q <= 32'b00000000000000000000000000000000 ;
        1337: q <= 32'b00000000000000000000000000000000 ;
        1338: q <= 32'b00000000000000000000000000000000 ;
        1339: q <= 32'b00000000000000000000000000000000 ;
        1340: q <= 32'b00000000000000000000000000000000 ;
        1341: q <= 32'b00000000000000000000000000000000 ;
        1342: q <= 32'b00000000000000000000000000000000 ;
        1343: q <= 32'b00000000000000000000000000000000 ;
        1344: q <= 32'b00000000000000000000000000000000 ;
        1345: q <= 32'b00000000000000000000000000000000 ;
        1346: q <= 32'b00000000000000000000000000000000 ;
        1347: q <= 32'b00000000000000000000000000000000 ;
        1348: q <= 32'b00000000000000000000000000000000 ;
        1349: q <= 32'b00000000000000000000000000000000 ;
        1350: q <= 32'b00000000000000000000000000000000 ;
        1351: q <= 32'b00000000000000000000000000000000 ;
        1352: q <= 32'b00000000000000000000000000000000 ;
        1353: q <= 32'b00000000000000000000000000000000 ;
        1354: q <= 32'b00000000000000000000000000000000 ;
        1355: q <= 32'b00000000000000000000000000000000 ;
        1356: q <= 32'b00000000000000000000000000000000 ;
        1357: q <= 32'b00000000000000000000000000000000 ;
        1358: q <= 32'b00000000000000000000000000000000 ;
        1359: q <= 32'b00000000000000000000000000000000 ;
        1360: q <= 32'b00000000000000000000000000000000 ;
        1361: q <= 32'b00000000000000000000000000000000 ;
        1362: q <= 32'b00000000000000000000000000000000 ;
        1363: q <= 32'b00000000000000000000000000000000 ;
        1364: q <= 32'b00000000000000000000000000000000 ;
        1365: q <= 32'b00000000000000000000000000000000 ;
        1366: q <= 32'b00000000000000000000000000000000 ;
        1367: q <= 32'b00000000000000000000000000000000 ;
        1368: q <= 32'b00000000000000000000000000000000 ;
        1369: q <= 32'b00000000000000000000000000000000 ;
        1370: q <= 32'b00000000000000000000000000000000 ;
        1371: q <= 32'b00000000000000000000000000000000 ;
        1372: q <= 32'b00000000000000000000000000000000 ;
        1373: q <= 32'b00000000000000000000000000000000 ;
        1374: q <= 32'b00000000000000000000000000000000 ;
        1375: q <= 32'b00000000000000000000000000000000 ;
        1376: q <= 32'b00000000000000000000000000000000 ;
        1377: q <= 32'b00000000000000000000000000000000 ;
        1378: q <= 32'b00000000000000000000000000000000 ;
        1379: q <= 32'b00000000000000000000000000000000 ;
        1380: q <= 32'b00000000000000000000000000000000 ;
        1381: q <= 32'b00000000000000000000000000000000 ;
        1382: q <= 32'b00000000000000000000000000000000 ;
        1383: q <= 32'b00000000000000000000000000000000 ;
        1384: q <= 32'b00000000000000000000000000000000 ;
        1385: q <= 32'b00000000000000000000000000000000 ;
        1386: q <= 32'b00000000000000000000000000000000 ;
        1387: q <= 32'b00000000000000000000000000000000 ;
        1388: q <= 32'b00000000000000000000000000000000 ;
        1389: q <= 32'b00000000000000000000000000000000 ;
        1390: q <= 32'b00000000000000000000000000000000 ;
        1391: q <= 32'b00000000000000000000000000000000 ;
        1392: q <= 32'b00000000000000000000000000000000 ;
        1393: q <= 32'b00000000000000000000000000000000 ;
        1394: q <= 32'b00000000000000000000000000000000 ;
        1395: q <= 32'b00000000000000000000000000000000 ;
        1396: q <= 32'b00000000000000000000000000000000 ;
        1397: q <= 32'b00000000000000000000000000000000 ;
        1398: q <= 32'b00000000000000000000000000000000 ;
        1399: q <= 32'b00000000000000000000000000000000 ;
        1400: q <= 32'b00000000000000000000000000000000 ;
        1401: q <= 32'b00000000000000000000000000000000 ;
        1402: q <= 32'b00000000000000000000000000000000 ;
        1403: q <= 32'b00000000000000000000000000000000 ;
        1404: q <= 32'b00000000000000000000000000000000 ;
        1405: q <= 32'b00000000000000000000000000000000 ;
        1406: q <= 32'b00000000000000000000000000000000 ;
        1407: q <= 32'b00000000000000000000000000000000 ;
        1408: q <= 32'b00000000000000000000000000000000 ;
        1409: q <= 32'b00000000000000000000000000000000 ;
        1410: q <= 32'b00000000000000000000000000000000 ;
        1411: q <= 32'b00000000000000000000000000000000 ;
        1412: q <= 32'b00000000000000000000000000000000 ;
        1413: q <= 32'b00000000000000000000000000000000 ;
        1414: q <= 32'b00000000000000000000000000000000 ;
        1415: q <= 32'b00000000000000000000000000000000 ;
        1416: q <= 32'b00000000000000000000000000000000 ;
        1417: q <= 32'b00000000000000000000000000000000 ;
        1418: q <= 32'b00000000000000000000000000000000 ;
        1419: q <= 32'b00000000000000000000000000000000 ;
        1420: q <= 32'b00000000000000000000000000000000 ;
        1421: q <= 32'b00000000000000000000000000000000 ;
        1422: q <= 32'b00000000000000000000000000000000 ;
        1423: q <= 32'b00000000000000000000000000000000 ;
        1424: q <= 32'b00000000000000000000000000000000 ;
        1425: q <= 32'b00000000000000000000000000000000 ;
        1426: q <= 32'b00000000000000000000000000000000 ;
        1427: q <= 32'b00000000000000000000000000000000 ;
        1428: q <= 32'b00000000000000000000000000000000 ;
        1429: q <= 32'b00000000000000000000000000000000 ;
        1430: q <= 32'b00000000000000000000000000000000 ;
        1431: q <= 32'b00000000000000000000000000000000 ;
        1432: q <= 32'b00000000000000000000000000000000 ;
        1433: q <= 32'b00000000000000000000000000000000 ;
        1434: q <= 32'b00000000000000000000000000000000 ;
        1435: q <= 32'b00000000000000000000000000000000 ;
        1436: q <= 32'b00000000000000000000000000000000 ;
        1437: q <= 32'b00000000000000000000000000000000 ;
        1438: q <= 32'b00000000000000000000000000000000 ;
        1439: q <= 32'b00000000000000000000000000000000 ;
        1440: q <= 32'b00000000000000000000000000000000 ;
        1441: q <= 32'b00000000000000000000000000000000 ;
        1442: q <= 32'b00000000000000000000000000000000 ;
        1443: q <= 32'b00000000000000000000000000000000 ;
        1444: q <= 32'b00000000000000000000000000000000 ;
        1445: q <= 32'b00000000000000000000000000000000 ;
        1446: q <= 32'b00000000000000000000000000000000 ;
        1447: q <= 32'b00000000000000000000000000000000 ;
        1448: q <= 32'b00000000000000000000000000000000 ;
        1449: q <= 32'b00000000000000000000000000000000 ;
        1450: q <= 32'b00000000000000000000000000000000 ;
        1451: q <= 32'b00000000000000000000000000000000 ;
        1452: q <= 32'b00000000000000000000000000000000 ;
        1453: q <= 32'b00000000000000000000000000000000 ;
        1454: q <= 32'b00000000000000000000000000000000 ;
        1455: q <= 32'b00000000000000000000000000000000 ;
        1456: q <= 32'b00000000000000000000000000000000 ;
        1457: q <= 32'b00000000000000000000000000000000 ;
        1458: q <= 32'b00000000000000000000000000000000 ;
        1459: q <= 32'b00000000000000000000000000000000 ;
        1460: q <= 32'b00000000000000000000000000000000 ;
        1461: q <= 32'b00000000000000000000000000000000 ;
        1462: q <= 32'b00000000000000000000000000000000 ;
        1463: q <= 32'b00000000000000000000000000000000 ;
        1464: q <= 32'b00000000000000000000000000000000 ;
        1465: q <= 32'b00000000000000000000000000000000 ;
        1466: q <= 32'b00000000000000000000000000000000 ;
        1467: q <= 32'b00000000000000000000000000000000 ;
        1468: q <= 32'b00000000000000000000000000000000 ;
        1469: q <= 32'b00000000000000000000000000000000 ;
        1470: q <= 32'b00000000000000000000000000000000 ;
        1471: q <= 32'b00000000000000000000000000000000 ;
        1472: q <= 32'b00000000000000000000000000000000 ;
        1473: q <= 32'b00000000000000000000000000000000 ;
        1474: q <= 32'b00000000000000000000000000000000 ;
        1475: q <= 32'b00000000000000000000000000000000 ;
        1476: q <= 32'b00000000000000000000000000000000 ;
        1477: q <= 32'b00000000000000000000000000000000 ;
        1478: q <= 32'b00000000000000000000000000000000 ;
        1479: q <= 32'b00000000000000000000000000000000 ;
        1480: q <= 32'b00000000000000000000000000000000 ;
        1481: q <= 32'b00000000000000000000000000000000 ;
        1482: q <= 32'b00000000000000000000000000000000 ;
        1483: q <= 32'b00000000000000000000000000000000 ;
        1484: q <= 32'b00000000000000000000000000000000 ;
        1485: q <= 32'b00000000000000000000000000000000 ;
        1486: q <= 32'b00000000000000000000000000000000 ;
        1487: q <= 32'b00000000000000000000000000000000 ;
        1488: q <= 32'b00000000000000000000000000000000 ;
        1489: q <= 32'b00000000000000000000000000000000 ;
        1490: q <= 32'b00000000000000000000000000000000 ;
        1491: q <= 32'b00000000000000000000000000000000 ;
        1492: q <= 32'b00000000000000000000000000000000 ;
        1493: q <= 32'b00000000000000000000000000000000 ;
        1494: q <= 32'b00000000000000000000000000000000 ;
        1495: q <= 32'b00000000000000000000000000000000 ;
        1496: q <= 32'b00000000000000000000000000000000 ;
        1497: q <= 32'b00000000000000000000000000000000 ;
        1498: q <= 32'b00000000000000000000000000000000 ;
        1499: q <= 32'b00000000000000000000000000000000 ;
        1500: q <= 32'b00000000000000000000000000000000 ;
        1501: q <= 32'b00000000000000000000000000000000 ;
        1502: q <= 32'b00000000000000000000000000000000 ;
        1503: q <= 32'b00000000000000000000000000000000 ;
        1504: q <= 32'b00000000000000000000000000000000 ;
        1505: q <= 32'b00000000000000000000000000000000 ;
        1506: q <= 32'b00000000000000000000000000000000 ;
        1507: q <= 32'b00000000000000000000000000000000 ;
        1508: q <= 32'b00000000000000000000000000000000 ;
        1509: q <= 32'b00000000000000000000000000000000 ;
        1510: q <= 32'b00000000000000000000000000000000 ;
        1511: q <= 32'b00000000000000000000000000000000 ;
        1512: q <= 32'b00000000000000000000000000000000 ;
        1513: q <= 32'b00000000000000000000000000000000 ;
        1514: q <= 32'b00000000000000000000000000000000 ;
        1515: q <= 32'b00000000000000000000000000000000 ;
        1516: q <= 32'b00000000000000000000000000000000 ;
        1517: q <= 32'b00000000000000000000000000000000 ;
        1518: q <= 32'b00000000000000000000000000000000 ;
        1519: q <= 32'b00000000000000000000000000000000 ;
        1520: q <= 32'b00000000000000000000000000000000 ;
        1521: q <= 32'b00000000000000000000000000000000 ;
        1522: q <= 32'b00000000000000000000000000000000 ;
        1523: q <= 32'b00000000000000000000000000000000 ;
        1524: q <= 32'b00000000000000000000000000000000 ;
        1525: q <= 32'b00000000000000000000000000000000 ;
        1526: q <= 32'b00000000000000000000000000000000 ;
        1527: q <= 32'b00000000000000000000000000000000 ;
        1528: q <= 32'b00000000000000000000000000000000 ;
        1529: q <= 32'b00000000000000000000000000000000 ;
        1530: q <= 32'b00000000000000000000000000000000 ;
        1531: q <= 32'b00000000000000000000000000000000 ;
        1532: q <= 32'b00000000000000000000000000000000 ;
        1533: q <= 32'b00000000000000000000000000000000 ;
        1534: q <= 32'b00000000000000000000000000000000 ;
        1535: q <= 32'b00000000000000000000000000000000 ;
        1536: q <= 32'b00000000000000000000000000000000 ;
        1537: q <= 32'b00000000000000000000000000000000 ;
        1538: q <= 32'b00000000000000000000000000000000 ;
        1539: q <= 32'b00000000000000000000000000000000 ;
        1540: q <= 32'b00000000000000000000000000000000 ;
        1541: q <= 32'b00000000000000000000000000000000 ;
        1542: q <= 32'b00000000000000000000000000000000 ;
        1543: q <= 32'b00000000000000000000000000000000 ;
        1544: q <= 32'b00000000000000000000000000000000 ;
        1545: q <= 32'b00000000000000000000000000000000 ;
        1546: q <= 32'b00000000000000000000000000000000 ;
        1547: q <= 32'b00000000000000000000000000000000 ;
        1548: q <= 32'b00000000000000000000000000000000 ;
        1549: q <= 32'b00000000000000000000000000000000 ;
        1550: q <= 32'b00000000000000000000000000000000 ;
        1551: q <= 32'b00000000000000000000000000000000 ;
        1552: q <= 32'b00000000000000000000000000000000 ;
        1553: q <= 32'b00000000000000000000000000000000 ;
        1554: q <= 32'b00000000000000000000000000000000 ;
        1555: q <= 32'b00000000000000000000000000000000 ;
        1556: q <= 32'b00000000000000000000000000000000 ;
        1557: q <= 32'b00000000000000000000000000000000 ;
        1558: q <= 32'b00000000000000000000000000000000 ;
        1559: q <= 32'b00000000000000000000000000000000 ;
        1560: q <= 32'b00000000000000000000000000000000 ;
        1561: q <= 32'b00000000000000000000000000000000 ;
        1562: q <= 32'b00000000000000000000000000000000 ;
        1563: q <= 32'b00000000000000000000000000000000 ;
        1564: q <= 32'b00000000000000000000000000000000 ;
        1565: q <= 32'b00000000000000000000000000000000 ;
        1566: q <= 32'b00000000000000000000000000000000 ;
        1567: q <= 32'b00000000000000000000000000000000 ;
        1568: q <= 32'b00000000000000000000000000000000 ;
        1569: q <= 32'b00000000000000000000000000000000 ;
        1570: q <= 32'b00000000000000000000000000000000 ;
        1571: q <= 32'b00000000000000000000000000000000 ;
        1572: q <= 32'b00000000000000000000000000000000 ;
        1573: q <= 32'b00000000000000000000000000000000 ;
        1574: q <= 32'b00000000000000000000000000000000 ;
        1575: q <= 32'b00000000000000000000000000000000 ;
        1576: q <= 32'b00000000000000000000000000000000 ;
        1577: q <= 32'b00000000000000000000000000000000 ;
        1578: q <= 32'b00000000000000000000000000000000 ;
        1579: q <= 32'b00000000000000000000000000000000 ;
        1580: q <= 32'b00000000000000000000000000000000 ;
        1581: q <= 32'b00000000000000000000000000000000 ;
        1582: q <= 32'b00000000000000000000000000000000 ;
        1583: q <= 32'b00000000000000000000000000000000 ;
        1584: q <= 32'b00000000000000000000000000000000 ;
        1585: q <= 32'b00000000000000000000000000000000 ;
        1586: q <= 32'b00000000000000000000000000000000 ;
        1587: q <= 32'b00000000000000000000000000000000 ;
        1588: q <= 32'b00000000000000000000000000000000 ;
        1589: q <= 32'b00000000000000000000000000000000 ;
        1590: q <= 32'b00000000000000000000000000000000 ;
        1591: q <= 32'b00000000000000000000000000000000 ;
        1592: q <= 32'b00000000000000000000000000000000 ;
        1593: q <= 32'b00000000000000000000000000000000 ;
        1594: q <= 32'b00000000000000000000000000000000 ;
        1595: q <= 32'b00000000000000000000000000000000 ;
        1596: q <= 32'b00000000000000000000000000000000 ;
        1597: q <= 32'b00000000000000000000000000000000 ;
        1598: q <= 32'b00000000000000000000000000000000 ;
        1599: q <= 32'b00000000000000000000000000000000 ;
        1600: q <= 32'b00000000000000000000000000000000 ;
        1601: q <= 32'b00000000000000000000000000000000 ;
        1602: q <= 32'b00000000000000000000000000000000 ;
        1603: q <= 32'b00000000000000000000000000000000 ;
        1604: q <= 32'b00000000000000000000000000000000 ;
        1605: q <= 32'b00000000000000000000000000000000 ;
        1606: q <= 32'b00000000000000000000000000000000 ;
        1607: q <= 32'b00000000000000000000000000000000 ;
        1608: q <= 32'b00000000000000000000000000000000 ;
        1609: q <= 32'b00000000000000000000000000000000 ;
        1610: q <= 32'b00000000000000000000000000000000 ;
        1611: q <= 32'b00000000000000000000000000000000 ;
        1612: q <= 32'b00000000000000000000000000000000 ;
        1613: q <= 32'b00000000000000000000000000000000 ;
        1614: q <= 32'b00000000000000000000000000000000 ;
        1615: q <= 32'b00000000000000000000000000000000 ;
        1616: q <= 32'b00000000000000000000000000000000 ;
        1617: q <= 32'b00000000000000000000000000000000 ;
        1618: q <= 32'b00000000000000000000000000000000 ;
        1619: q <= 32'b00000000000000000000000000000000 ;
        1620: q <= 32'b00000000000000000000000000000000 ;
        1621: q <= 32'b00000000000000000000000000000000 ;
        1622: q <= 32'b00000000000000000000000000000000 ;
        1623: q <= 32'b00000000000000000000000000000000 ;
        1624: q <= 32'b00000000000000000000000000000000 ;
        1625: q <= 32'b00000000000000000000000000000000 ;
        1626: q <= 32'b00000000000000000000000000000000 ;
        1627: q <= 32'b00000000000000000000000000000000 ;
        1628: q <= 32'b00000000000000000000000000000000 ;
        1629: q <= 32'b00000000000000000000000000000000 ;
        1630: q <= 32'b00000000000000000000000000000000 ;
        1631: q <= 32'b00000000000000000000000000000000 ;
        1632: q <= 32'b00000000000000000000000000000000 ;
        1633: q <= 32'b00000000000000000000000000000000 ;
        1634: q <= 32'b00000000000000000000000000000000 ;
        1635: q <= 32'b00000000000000000000000000000000 ;
        1636: q <= 32'b00000000000000000000000000000000 ;
        1637: q <= 32'b00000000000000000000000000000000 ;
        1638: q <= 32'b00000000000000000000000000000000 ;
        1639: q <= 32'b00000000000000000000000000000000 ;
        1640: q <= 32'b00000000000000000000000000000000 ;
        1641: q <= 32'b00000000000000000000000000000000 ;
        1642: q <= 32'b00000000000000000000000000000000 ;
        1643: q <= 32'b00000000000000000000000000000000 ;
        1644: q <= 32'b00000000000000000000000000000000 ;
        1645: q <= 32'b00000000000000000000000000000000 ;
        1646: q <= 32'b00000000000000000000000000000000 ;
        1647: q <= 32'b00000000000000000000000000000000 ;
        1648: q <= 32'b00000000000000000000000000000000 ;
        1649: q <= 32'b00000000000000000000000000000000 ;
        1650: q <= 32'b00000000000000000000000000000000 ;
        1651: q <= 32'b00000000000000000000000000000000 ;
        1652: q <= 32'b00000000000000000000000000000000 ;
        1653: q <= 32'b00000000000000000000000000000000 ;
        1654: q <= 32'b00000000000000000000000000000000 ;
        1655: q <= 32'b00000000000000000000000000000000 ;
        1656: q <= 32'b00000000000000000000000000000000 ;
        1657: q <= 32'b00000000000000000000000000000000 ;
        1658: q <= 32'b00000000000000000000000000000000 ;
        1659: q <= 32'b00000000000000000000000000000000 ;
        1660: q <= 32'b00000000000000000000000000000000 ;
        1661: q <= 32'b00000000000000000000000000000000 ;
        1662: q <= 32'b00000000000000000000000000000000 ;
        1663: q <= 32'b00000000000000000000000000000000 ;
        1664: q <= 32'b00000000000000000000000000000000 ;
        1665: q <= 32'b00000000000000000000000000000000 ;
        1666: q <= 32'b00000000000000000000000000000000 ;
        1667: q <= 32'b00000000000000000000000000000000 ;
        1668: q <= 32'b00000000000000000000000000000000 ;
        1669: q <= 32'b00000000000000000000000000000000 ;
        1670: q <= 32'b00000000000000000000000000000000 ;
        1671: q <= 32'b00000000000000000000000000000000 ;
        1672: q <= 32'b00000000000000000000000000000000 ;
        1673: q <= 32'b00000000000000000000000000000000 ;
        1674: q <= 32'b00000000000000000000000000000000 ;
        1675: q <= 32'b00000000000000000000000000000000 ;
        1676: q <= 32'b00000000000000000000000000000000 ;
        1677: q <= 32'b00000000000000000000000000000000 ;
        1678: q <= 32'b00000000000000000000000000000000 ;
        1679: q <= 32'b00000000000000000000000000000000 ;
        1680: q <= 32'b00000000000000000000000000000000 ;
        1681: q <= 32'b00000000000000000000000000000000 ;
        1682: q <= 32'b00000000000000000000000000000000 ;
        1683: q <= 32'b00000000000000000000000000000000 ;
        1684: q <= 32'b00000000000000000000000000000000 ;
        1685: q <= 32'b00000000000000000000000000000000 ;
        1686: q <= 32'b00000000000000000000000000000000 ;
        1687: q <= 32'b00000000000000000000000000000000 ;
        1688: q <= 32'b00000000000000000000000000000000 ;
        1689: q <= 32'b00000000000000000000000000000000 ;
        1690: q <= 32'b00000000000000000000000000000000 ;
        1691: q <= 32'b00000000000000000000000000000000 ;
        1692: q <= 32'b00000000000000000000000000000000 ;
        1693: q <= 32'b00000000000000000000000000000000 ;
        1694: q <= 32'b00000000000000000000000000000000 ;
        1695: q <= 32'b00000000000000000000000000000000 ;
        1696: q <= 32'b00000000000000000000000000000000 ;
        1697: q <= 32'b00000000000000000000000000000000 ;
        1698: q <= 32'b00000000000000000000000000000000 ;
        1699: q <= 32'b00000000000000000000000000000000 ;
        1700: q <= 32'b00000000000000000000000000000000 ;
        1701: q <= 32'b00000000000000000000000000000000 ;
        1702: q <= 32'b00000000000000000000000000000000 ;
        1703: q <= 32'b00000000000000000000000000000000 ;
        1704: q <= 32'b00000000000000000000000000000000 ;
        1705: q <= 32'b00000000000000000000000000000000 ;
        1706: q <= 32'b00000000000000000000000000000000 ;
        1707: q <= 32'b00000000000000000000000000000000 ;
        1708: q <= 32'b00000000000000000000000000000000 ;
        1709: q <= 32'b00000000000000000000000000000000 ;
        1710: q <= 32'b00000000000000000000000000000000 ;
        1711: q <= 32'b00000000000000000000000000000000 ;
        1712: q <= 32'b00000000000000000000000000000000 ;
        1713: q <= 32'b00000000000000000000000000000000 ;
        1714: q <= 32'b00000000000000000000000000000000 ;
        1715: q <= 32'b00000000000000000000000000000000 ;
        1716: q <= 32'b00000000000000000000000000000000 ;
        1717: q <= 32'b00000000000000000000000000000000 ;
        1718: q <= 32'b00000000000000000000000000000000 ;
        1719: q <= 32'b00000000000000000000000000000000 ;
        1720: q <= 32'b00000000000000000000000000000000 ;
        1721: q <= 32'b00000000000000000000000000000000 ;
        1722: q <= 32'b00000000000000000000000000000000 ;
        1723: q <= 32'b00000000000000000000000000000000 ;
        1724: q <= 32'b00000000000000000000000000000000 ;
        1725: q <= 32'b00000000000000000000000000000000 ;
        1726: q <= 32'b00000000000000000000000000000000 ;
        1727: q <= 32'b00000000000000000000000000000000 ;
        1728: q <= 32'b00000000000000000000000000000000 ;
        1729: q <= 32'b00000000000000000000000000000000 ;
        1730: q <= 32'b00000000000000000000000000000000 ;
        1731: q <= 32'b00000000000000000000000000000000 ;
        1732: q <= 32'b00000000000000000000000000000000 ;
        1733: q <= 32'b00000000000000000000000000000000 ;
        1734: q <= 32'b00000000000000000000000000000000 ;
        1735: q <= 32'b00000000000000000000000000000000 ;
        1736: q <= 32'b00000000000000000000000000000000 ;
        1737: q <= 32'b00000000000000000000000000000000 ;
        1738: q <= 32'b00000000000000000000000000000000 ;
        1739: q <= 32'b00000000000000000000000000000000 ;
        1740: q <= 32'b00000000000000000000000000000000 ;
        1741: q <= 32'b00000000000000000000000000000000 ;
        1742: q <= 32'b00000000000000000000000000000000 ;
        1743: q <= 32'b00000000000000000000000000000000 ;
        1744: q <= 32'b00000000000000000000000000000000 ;
        1745: q <= 32'b00000000000000000000000000000000 ;
        1746: q <= 32'b00000000000000000000000000000000 ;
        1747: q <= 32'b00000000000000000000000000000000 ;
        1748: q <= 32'b00000000000000000000000000000000 ;
        1749: q <= 32'b00000000000000000000000000000000 ;
        1750: q <= 32'b00000000000000000000000000000000 ;
        1751: q <= 32'b00000000000000000000000000000000 ;
        1752: q <= 32'b00000000000000000000000000000000 ;
        1753: q <= 32'b00000000000000000000000000000000 ;
        1754: q <= 32'b00000000000000000000000000000000 ;
        1755: q <= 32'b00000000000000000000000000000000 ;
        1756: q <= 32'b00000000000000000000000000000000 ;
        1757: q <= 32'b00000000000000000000000000000000 ;
        1758: q <= 32'b00000000000000000000000000000000 ;
        1759: q <= 32'b00000000000000000000000000000000 ;
        1760: q <= 32'b00000000000000000000000000000000 ;
        1761: q <= 32'b00000000000000000000000000000000 ;
        1762: q <= 32'b00000000000000000000000000000000 ;
        1763: q <= 32'b00000000000000000000000000000000 ;
        1764: q <= 32'b00000000000000000000000000000000 ;
        1765: q <= 32'b00000000000000000000000000000000 ;
        1766: q <= 32'b00000000000000000000000000000000 ;
        1767: q <= 32'b00000000000000000000000000000000 ;
        1768: q <= 32'b00000000000000000000000000000000 ;
        1769: q <= 32'b00000000000000000000000000000000 ;
        1770: q <= 32'b00000000000000000000000000000000 ;
        1771: q <= 32'b00000000000000000000000000000000 ;
        1772: q <= 32'b00000000000000000000000000000000 ;
        1773: q <= 32'b00000000000000000000000000000000 ;
        1774: q <= 32'b00000000000000000000000000000000 ;
        1775: q <= 32'b00000000000000000000000000000000 ;
        1776: q <= 32'b00000000000000000000000000000000 ;
        1777: q <= 32'b00000000000000000000000000000000 ;
        1778: q <= 32'b00000000000000000000000000000000 ;
        1779: q <= 32'b00000000000000000000000000000000 ;
        1780: q <= 32'b00000000000000000000000000000000 ;
        1781: q <= 32'b00000000000000000000000000000000 ;
        1782: q <= 32'b00000000000000000000000000000000 ;
        1783: q <= 32'b00000000000000000000000000000000 ;
        1784: q <= 32'b00000000000000000000000000000000 ;
        1785: q <= 32'b00000000000000000000000000000000 ;
        1786: q <= 32'b00000000000000000000000000000000 ;
        1787: q <= 32'b00000000000000000000000000000000 ;
        1788: q <= 32'b00000000000000000000000000000000 ;
        1789: q <= 32'b00000000000000000000000000000000 ;
        1790: q <= 32'b00000000000000000000000000000000 ;
        1791: q <= 32'b00000000000000000000000000000000 ;
        1792: q <= 32'b00000000000000000000000000000000 ;
        1793: q <= 32'b00000000000000000000000000000000 ;
        1794: q <= 32'b00000000000000000000000000000000 ;
        1795: q <= 32'b00000000000000000000000000000000 ;
        1796: q <= 32'b00000000000000000000000000000000 ;
        1797: q <= 32'b00000000000000000000000000000000 ;
        1798: q <= 32'b00000000000000000000000000000000 ;
        1799: q <= 32'b00000000000000000000000000000000 ;
        1800: q <= 32'b00000000000000000000000000000000 ;
        1801: q <= 32'b00000000000000000000000000000000 ;
        1802: q <= 32'b00000000000000000000000000000000 ;
        1803: q <= 32'b00000000000000000000000000000000 ;
        1804: q <= 32'b00000000000000000000000000000000 ;
        1805: q <= 32'b00000000000000000000000000000000 ;
        1806: q <= 32'b00000000000000000000000000000000 ;
        1807: q <= 32'b00000000000000000000000000000000 ;
        1808: q <= 32'b00000000000000000000000000000000 ;
        1809: q <= 32'b00000000000000000000000000000000 ;
        1810: q <= 32'b00000000000000000000000000000000 ;
        1811: q <= 32'b00000000000000000000000000000000 ;
        1812: q <= 32'b00000000000000000000000000000000 ;
        1813: q <= 32'b00000000000000000000000000000000 ;
        1814: q <= 32'b00000000000000000000000000000000 ;
        1815: q <= 32'b00000000000000000000000000000000 ;
        1816: q <= 32'b00000000000000000000000000000000 ;
        1817: q <= 32'b00000000000000000000000000000000 ;
        1818: q <= 32'b00000000000000000000000000000000 ;
        1819: q <= 32'b00000000000000000000000000000000 ;
        1820: q <= 32'b00000000000000000000000000000000 ;
        1821: q <= 32'b00000000000000000000000000000000 ;
        1822: q <= 32'b00000000000000000000000000000000 ;
        1823: q <= 32'b00000000000000000000000000000000 ;
        1824: q <= 32'b00000000000000000000000000000000 ;
        1825: q <= 32'b00000000000000000000000000000000 ;
        1826: q <= 32'b00000000000000000000000000000000 ;
        1827: q <= 32'b00000000000000000000000000000000 ;
        1828: q <= 32'b00000000000000000000000000000000 ;
        1829: q <= 32'b00000000000000000000000000000000 ;
        1830: q <= 32'b00000000000000000000000000000000 ;
        1831: q <= 32'b00000000000000000000000000000000 ;
        1832: q <= 32'b00000000000000000000000000000000 ;
        1833: q <= 32'b00000000000000000000000000000000 ;
        1834: q <= 32'b00000000000000000000000000000000 ;
        1835: q <= 32'b00000000000000000000000000000000 ;
        1836: q <= 32'b00000000000000000000000000000000 ;
        1837: q <= 32'b00000000000000000000000000000000 ;
        1838: q <= 32'b00000000000000000000000000000000 ;
        1839: q <= 32'b00000000000000000000000000000000 ;
        1840: q <= 32'b00000000000000000000000000000000 ;
        1841: q <= 32'b00000000000000000000000000000000 ;
        1842: q <= 32'b00000000000000000000000000000000 ;
        1843: q <= 32'b00000000000000000000000000000000 ;
        1844: q <= 32'b00000000000000000000000000000000 ;
        1845: q <= 32'b00000000000000000000000000000000 ;
        1846: q <= 32'b00000000000000000000000000000000 ;
        1847: q <= 32'b00000000000000000000000000000000 ;
        1848: q <= 32'b00000000000000000000000000000000 ;
        1849: q <= 32'b00000000000000000000000000000000 ;
        1850: q <= 32'b00000000000000000000000000000000 ;
        1851: q <= 32'b00000000000000000000000000000000 ;
        1852: q <= 32'b00000000000000000000000000000000 ;
        1853: q <= 32'b00000000000000000000000000000000 ;
        1854: q <= 32'b00000000000000000000000000000000 ;
        1855: q <= 32'b00000000000000000000000000000000 ;
        1856: q <= 32'b00000000000000000000000000000000 ;
        1857: q <= 32'b00000000000000000000000000000000 ;
        1858: q <= 32'b00000000000000000000000000000000 ;
        1859: q <= 32'b00000000000000000000000000000000 ;
        1860: q <= 32'b00000000000000000000000000000000 ;
        1861: q <= 32'b00000000000000000000000000000000 ;
        1862: q <= 32'b00000000000000000000000000000000 ;
        1863: q <= 32'b00000000000000000000000000000000 ;
        1864: q <= 32'b00000000000000000000000000000000 ;
        1865: q <= 32'b00000000000000000000000000000000 ;
        1866: q <= 32'b00000000000000000000000000000000 ;
        1867: q <= 32'b00000000000000000000000000000000 ;
        1868: q <= 32'b00000000000000000000000000000000 ;
        1869: q <= 32'b00000000000000000000000000000000 ;
        1870: q <= 32'b00000000000000000000000000000000 ;
        1871: q <= 32'b00000000000000000000000000000000 ;
        1872: q <= 32'b00000000000000000000000000000000 ;
        1873: q <= 32'b00000000000000000000000000000000 ;
        1874: q <= 32'b00000000000000000000000000000000 ;
        1875: q <= 32'b00000000000000000000000000000000 ;
        1876: q <= 32'b00000000000000000000000000000000 ;
        1877: q <= 32'b00000000000000000000000000000000 ;
        1878: q <= 32'b00000000000000000000000000000000 ;
        1879: q <= 32'b00000000000000000000000000000000 ;
        1880: q <= 32'b00000000000000000000000000000000 ;
        1881: q <= 32'b00000000000000000000000000000000 ;
        1882: q <= 32'b00000000000000000000000000000000 ;
        1883: q <= 32'b00000000000000000000000000000000 ;
        1884: q <= 32'b00000000000000000000000000000000 ;
        1885: q <= 32'b00000000000000000000000000000000 ;
        1886: q <= 32'b00000000000000000000000000000000 ;
        1887: q <= 32'b00000000000000000000000000000000 ;
        1888: q <= 32'b00000000000000000000000000000000 ;
        1889: q <= 32'b00000000000000000000000000000000 ;
        1890: q <= 32'b00000000000000000000000000000000 ;
        1891: q <= 32'b00000000000000000000000000000000 ;
        1892: q <= 32'b00000000000000000000000000000000 ;
        1893: q <= 32'b00000000000000000000000000000000 ;
        1894: q <= 32'b00000000000000000000000000000000 ;
        1895: q <= 32'b00000000000000000000000000000000 ;
        1896: q <= 32'b00000000000000000000000000000000 ;
        1897: q <= 32'b00000000000000000000000000000000 ;
        1898: q <= 32'b00000000000000000000000000000000 ;
        1899: q <= 32'b00000000000000000000000000000000 ;
        1900: q <= 32'b00000000000000000000000000000000 ;
        1901: q <= 32'b00000000000000000000000000000000 ;
        1902: q <= 32'b00000000000000000000000000000000 ;
        1903: q <= 32'b00000000000000000000000000000000 ;
        1904: q <= 32'b00000000000000000000000000000000 ;
        1905: q <= 32'b00000000000000000000000000000000 ;
        1906: q <= 32'b00000000000000000000000000000000 ;
        1907: q <= 32'b00000000000000000000000000000000 ;
        1908: q <= 32'b00000000000000000000000000000000 ;
        1909: q <= 32'b00000000000000000000000000000000 ;
        1910: q <= 32'b00000000000000000000000000000000 ;
        1911: q <= 32'b00000000000000000000000000000000 ;
        1912: q <= 32'b00000000000000000000000000000000 ;
        1913: q <= 32'b00000000000000000000000000000000 ;
        1914: q <= 32'b00000000000000000000000000000000 ;
        1915: q <= 32'b00000000000000000000000000000000 ;
        1916: q <= 32'b00000000000000000000000000000000 ;
        1917: q <= 32'b00000000000000000000000000000000 ;
        1918: q <= 32'b00000000000000000000000000000000 ;
        1919: q <= 32'b00000000000000000000000000000000 ;
        1920: q <= 32'b00000000000000000000000000000000 ;
        1921: q <= 32'b00000000000000000000000000000000 ;
        1922: q <= 32'b00000000000000000000000000000000 ;
        1923: q <= 32'b00000000000000000000000000000000 ;
        1924: q <= 32'b00000000000000000000000000000000 ;
        1925: q <= 32'b00000000000000000000000000000000 ;
        1926: q <= 32'b00000000000000000000000000000000 ;
        1927: q <= 32'b00000000000000000000000000000000 ;
        1928: q <= 32'b00000000000000000000000000000000 ;
        1929: q <= 32'b00000000000000000000000000000000 ;
        1930: q <= 32'b00000000000000000000000000000000 ;
        1931: q <= 32'b00000000000000000000000000000000 ;
        1932: q <= 32'b00000000000000000000000000000000 ;
        1933: q <= 32'b00000000000000000000000000000000 ;
        1934: q <= 32'b00000000000000000000000000000000 ;
        1935: q <= 32'b00000000000000000000000000000000 ;
        1936: q <= 32'b00000000000000000000000000000000 ;
        1937: q <= 32'b00000000000000000000000000000000 ;
        1938: q <= 32'b00000000000000000000000000000000 ;
        1939: q <= 32'b00000000000000000000000000000000 ;
        1940: q <= 32'b00000000000000000000000000000000 ;
        1941: q <= 32'b00000000000000000000000000000000 ;
        1942: q <= 32'b00000000000000000000000000000000 ;
        1943: q <= 32'b00000000000000000000000000000000 ;
        1944: q <= 32'b00000000000000000000000000000000 ;
        1945: q <= 32'b00000000000000000000000000000000 ;
        1946: q <= 32'b00000000000000000000000000000000 ;
        1947: q <= 32'b00000000000000000000000000000000 ;
        1948: q <= 32'b00000000000000000000000000000000 ;
        1949: q <= 32'b00000000000000000000000000000000 ;
        1950: q <= 32'b00000000000000000000000000000000 ;
        1951: q <= 32'b00000000000000000000000000000000 ;
        1952: q <= 32'b00000000000000000000000000000000 ;
        1953: q <= 32'b00000000000000000000000000000000 ;
        1954: q <= 32'b00000000000000000000000000000000 ;
        1955: q <= 32'b00000000000000000000000000000000 ;
        1956: q <= 32'b00000000000000000000000000000000 ;
        1957: q <= 32'b00000000000000000000000000000000 ;
        1958: q <= 32'b00000000000000000000000000000000 ;
        1959: q <= 32'b00000000000000000000000000000000 ;
        1960: q <= 32'b00000000000000000000000000000000 ;
        1961: q <= 32'b00000000000000000000000000000000 ;
        1962: q <= 32'b00000000000000000000000000000000 ;
        1963: q <= 32'b00000000000000000000000000000000 ;
        1964: q <= 32'b00000000000000000000000000000000 ;
        1965: q <= 32'b00000000000000000000000000000000 ;
        1966: q <= 32'b00000000000000000000000000000000 ;
        1967: q <= 32'b00000000000000000000000000000000 ;
        1968: q <= 32'b00000000000000000000000000000000 ;
        1969: q <= 32'b00000000000000000000000000000000 ;
        1970: q <= 32'b00000000000000000000000000000000 ;
        1971: q <= 32'b00000000000000000000000000000000 ;
        1972: q <= 32'b00000000000000000000000000000000 ;
        1973: q <= 32'b00000000000000000000000000000000 ;
        1974: q <= 32'b00000000000000000000000000000000 ;
        1975: q <= 32'b00000000000000000000000000000000 ;
        1976: q <= 32'b00000000000000000000000000000000 ;
        1977: q <= 32'b00000000000000000000000000000000 ;
        1978: q <= 32'b00000000000000000000000000000000 ;
        1979: q <= 32'b00000000000000000000000000000000 ;
        1980: q <= 32'b00000000000000000000000000000000 ;
        1981: q <= 32'b00000000000000000000000000000000 ;
        1982: q <= 32'b00000000000000000000000000000000 ;
        1983: q <= 32'b00000000000000000000000000000000 ;
        1984: q <= 32'b00000000000000000000000000000000 ;
        1985: q <= 32'b00000000000000000000000000000000 ;
        1986: q <= 32'b00000000000000000000000000000000 ;
        1987: q <= 32'b00000000000000000000000000000000 ;
        1988: q <= 32'b00000000000000000000000000000000 ;
        1989: q <= 32'b00000000000000000000000000000000 ;
        1990: q <= 32'b00000000000000000000000000000000 ;
        1991: q <= 32'b00000000000000000000000000000000 ;
        1992: q <= 32'b00000000000000000000000000000000 ;
        1993: q <= 32'b00000000000000000000000000000000 ;
        1994: q <= 32'b00000000000000000000000000000000 ;
        1995: q <= 32'b00000000000000000000000000000000 ;
        1996: q <= 32'b00000000000000000000000000000000 ;
        1997: q <= 32'b00000000000000000000000000000000 ;
        1998: q <= 32'b00000000000000000000000000000000 ;
        1999: q <= 32'b00000000000000000000000000000000 ;
        2000: q <= 32'b00000000000000000000000000000000 ;
        2001: q <= 32'b00000000000000000000000000000000 ;
        2002: q <= 32'b00000000000000000000000000000000 ;
        2003: q <= 32'b00000000000000000000000000000000 ;
        2004: q <= 32'b00000000000000000000000000000000 ;
        2005: q <= 32'b00000000000000000000000000000000 ;
        2006: q <= 32'b00000000000000000000000000000000 ;
        2007: q <= 32'b00000000000000000000000000000000 ;
        2008: q <= 32'b00000000000000000000000000000000 ;
        2009: q <= 32'b00000000000000000000000000000000 ;
        2010: q <= 32'b00000000000000000000000000000000 ;
        2011: q <= 32'b00000000000000000000000000000000 ;
        2012: q <= 32'b00000000000000000000000000000000 ;
        2013: q <= 32'b00000000000000000000000000000000 ;
        2014: q <= 32'b00000000000000000000000000000000 ;
        2015: q <= 32'b00000000000000000000000000000000 ;
        2016: q <= 32'b00000000000000000000000000000000 ;
        2017: q <= 32'b00000000000000000000000000000000 ;
        2018: q <= 32'b00000000000000000000000000000000 ;
        2019: q <= 32'b00000000000000000000000000000000 ;
        2020: q <= 32'b00000000000000000000000000000000 ;
        2021: q <= 32'b00000000000000000000000000000000 ;
        2022: q <= 32'b00000000000000000000000000000000 ;
        2023: q <= 32'b00000000000000000000000000000000 ;
        2024: q <= 32'b00000000000000000000000000000000 ;
        2025: q <= 32'b00000000000000000000000000000000 ;
        2026: q <= 32'b00000000000000000000000000000000 ;
        2027: q <= 32'b00000000000000000000000000000000 ;
        2028: q <= 32'b00000000000000000000000000000000 ;
        2029: q <= 32'b00000000000000000000000000000000 ;
        2030: q <= 32'b00000000000000000000000000000000 ;
        2031: q <= 32'b00000000000000000000000000000000 ;
        2032: q <= 32'b00000000000000000000000000000000 ;
        2033: q <= 32'b00000000000000000000000000000000 ;
        2034: q <= 32'b00000000000000000000000000000000 ;
        2035: q <= 32'b00000000000000000000000000000000 ;
        2036: q <= 32'b00000000000000000000000000000000 ;
        2037: q <= 32'b00000000000000000000000000000000 ;
        2038: q <= 32'b00000000000000000000000000000000 ;
        2039: q <= 32'b00000000000000000000000000000000 ;
        2040: q <= 32'b00000000000000000000000000000000 ;
        2041: q <= 32'b00000000000000000000000000000000 ;
        2042: q <= 32'b00000000000000000000000000000000 ;
        2043: q <= 32'b00000000000000000000000000000000 ;
        2044: q <= 32'b00000000000000000000000000000000 ;
        2045: q <= 32'b00000000000000000000000000000000 ;
        2046: q <= 32'b00000000000000000000000000000000 ;
        2047: q <= 32'b00000000000000000000000000000000 ;
        default: q <= 32'b00000000000000000000000000000000;
    endcase
end

endmodule
