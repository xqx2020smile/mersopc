module mem_rom_weight_out_01 (clock, address, q) ;
parameter DATA_WIDTH =  32;
input clock;
input [9:0] address;
output [DATA_WIDTH-1:0] q;
reg    [DATA_WIDTH-1:0] q;
always@(posedge clock) begin 
    case(address)
        0: q <= 32'b00111110000111111100101011101011 ;
        1: q <= 32'b10111110111011100110111010101101 ;
        2: q <= 32'b00111111000010000111001000001001 ;
        3: q <= 32'b00111101001010001101011101000010 ;
        4: q <= 32'b00111110100010100011100001110001 ;
        5: q <= 32'b00111110101111001010001111010110 ;
        6: q <= 32'b10111110100010111010001111000101 ;
        7: q <= 32'b10111110100111000001011000110111 ;
        8: q <= 32'b00111110011001110101111101100101 ;
        9: q <= 32'b10111111000001100101000111001101 ;
        10: q <= 32'b10111111001011001010010101001010 ;
        11: q <= 32'b00111101100000001011000011101011 ;
        12: q <= 32'b00111110001010011000100011100100 ;
        13: q <= 32'b10111110100011001111010011011110 ;
        14: q <= 32'b10111110110101001101101001000010 ;
        15: q <= 32'b10111110000000101111001101001110 ;
        16: q <= 32'b10111110000001001101010011000011 ;
        17: q <= 32'b00111110100101110111101011010001 ;
        18: q <= 32'b10111110110011111110110010110110 ;
        19: q <= 32'b00111110100010101010101011001110 ;
        20: q <= 32'b10111111001011000111011111111101 ;
        21: q <= 32'b00111101011011000111101001101100 ;
        22: q <= 32'b10111110000100100101111101111001 ;
        23: q <= 32'b00111110001010001111010110111001 ;
        24: q <= 32'b00111110001111011110101111010010 ;
        25: q <= 32'b10111110010011111011101001010110 ;
        26: q <= 32'b10111110110011111101010010111110 ;
        27: q <= 32'b00111110100101011100001100100001 ;
        28: q <= 32'b00111101100110001000001010101001 ;
        29: q <= 32'b10111110100100001100110101000010 ;
        30: q <= 32'b00111101111011011001011011101110 ;
        31: q <= 32'b10111101101110110010000111001111 ;
        32: q <= 32'b10111110010100110011001011111010 ;
        33: q <= 32'b10111110011110011110011001110110 ;
        34: q <= 32'b00111111001011000111011111001000 ;
        35: q <= 32'b00111111000010010111100011101100 ;
        36: q <= 32'b00111110100011110101001011011100 ;
        37: q <= 32'b00111110000010011110010101100110 ;
        38: q <= 32'b00111101010000000001010100110011 ;
        39: q <= 32'b00111110111101010111110100011100 ;
        40: q <= 32'b10111110010010011110110000010000 ;
        41: q <= 32'b10111111000101010101100000011000 ;
        42: q <= 32'b00111110011010110110011010010110 ;
        43: q <= 32'b00111111000001100010111000110100 ;
        44: q <= 32'b00111101111001011000101111100010 ;
        45: q <= 32'b00111101001110000111100001110110 ;
        46: q <= 32'b00111101110100110111110100100000 ;
        47: q <= 32'b00111101110001010010100101110101 ;
        48: q <= 32'b00111110010110001000111010111001 ;
        49: q <= 32'b10111010111111011011101101111100 ;
        50: q <= 32'b10111110011011010011010000111011 ;
        51: q <= 32'b10111101010001001110101111110011 ;
        52: q <= 32'b10111110001010110010101110011010 ;
        53: q <= 32'b10111110000001110001100100011111 ;
        54: q <= 32'b00111110010100111000111110000011 ;
        55: q <= 32'b00111110100000011101001011101111 ;
        56: q <= 32'b00111011101001100101011011100101 ;
        57: q <= 32'b10111110100000110111110111011100 ;
        58: q <= 32'b00111110100001001001011111000110 ;
        59: q <= 32'b10111110100101110011000000101010 ;
        60: q <= 32'b00000000000000000000000000000000 ;
        61: q <= 32'b00000000000000000000000000000000 ;
        62: q <= 32'b00000000000000000000000000000000 ;
        63: q <= 32'b00000000000000000000000000000000 ;
        64: q <= 32'b00111101001100110110010010011001 ;
        65: q <= 32'b00111110000110100000011101100110 ;
        66: q <= 32'b00111111000111001010011110000110 ;
        67: q <= 32'b10111101110011111101110100010001 ;
        68: q <= 32'b00111101011111100000100000001111 ;
        69: q <= 32'b00111110100000101011100001010110 ;
        70: q <= 32'b10111101010010111001111110001100 ;
        71: q <= 32'b10111110011110111111111011011100 ;
        72: q <= 32'b10111110111101010001111000011110 ;
        73: q <= 32'b10111101101111100100101001100010 ;
        74: q <= 32'b00111101100011010110010100001011 ;
        75: q <= 32'b10111111010010101001110110011111 ;
        76: q <= 32'b00111101010011011110010101011000 ;
        77: q <= 32'b10111110001101100110110110101001 ;
        78: q <= 32'b10111111000100001101110111100000 ;
        79: q <= 32'b10111110101000100111011011111011 ;
        80: q <= 32'b10111110000111011010000100100110 ;
        81: q <= 32'b00111111000001010011011100000111 ;
        82: q <= 32'b00111110101111010111101111011101 ;
        83: q <= 32'b10111101101100001111011111101010 ;
        84: q <= 32'b00111101110011100001110010100111 ;
        85: q <= 32'b10111101100010011000110110100111 ;
        86: q <= 32'b00111110110000011000111000111011 ;
        87: q <= 32'b00111110010000110101000100110010 ;
        88: q <= 32'b10111111001110101111101001000100 ;
        89: q <= 32'b00111100110110111110111000011010 ;
        90: q <= 32'b00111110111101011110100000000111 ;
        91: q <= 32'b00111110001000011110010011000000 ;
        92: q <= 32'b00111110011011001111001000100101 ;
        93: q <= 32'b10111110010011110100001000101000 ;
        94: q <= 32'b00111110011001010101111110111101 ;
        95: q <= 32'b10111101110100110110001010011110 ;
        96: q <= 32'b00111111000000100101111111101001 ;
        97: q <= 32'b10111101111110111111110111111101 ;
        98: q <= 32'b00111110111010011000110011000000 ;
        99: q <= 32'b00111110011011011011101000100100 ;
        100: q <= 32'b00111101100011011001011100000011 ;
        101: q <= 32'b00111110010110101101011101100100 ;
        102: q <= 32'b10111111010010010110010001010010 ;
        103: q <= 32'b00111101100000000001010001000010 ;
        104: q <= 32'b10111101101001110101001010011100 ;
        105: q <= 32'b00111110011001111001110110110100 ;
        106: q <= 32'b00111110100101010111111110111110 ;
        107: q <= 32'b10111110010111110011111111001001 ;
        108: q <= 32'b00111110000111001011010101011111 ;
        109: q <= 32'b10111101101000011001001000100101 ;
        110: q <= 32'b10111100010100011100011111110010 ;
        111: q <= 32'b00111101111110101001010110011010 ;
        112: q <= 32'b00111101110010011001101000001001 ;
        113: q <= 32'b00111100110001111100100101111111 ;
        114: q <= 32'b10111101110000010111111110001110 ;
        115: q <= 32'b00111100100101111001111110101001 ;
        116: q <= 32'b00111101011100011110000111110000 ;
        117: q <= 32'b10111110101001000101011110011101 ;
        118: q <= 32'b00111011100010110010100000110100 ;
        119: q <= 32'b10111011101110101011110011000001 ;
        120: q <= 32'b00111111001000011001010000000110 ;
        121: q <= 32'b10111110010001001010111110111110 ;
        122: q <= 32'b00111110111110010000111110110101 ;
        123: q <= 32'b10111110010110000101011110000010 ;
        124: q <= 32'b00000000000000000000000000000000 ;
        125: q <= 32'b00000000000000000000000000000000 ;
        126: q <= 32'b00000000000000000000000000000000 ;
        127: q <= 32'b00000000000000000000000000000000 ;
        128: q <= 32'b00111110100111000110011001011011 ;
        129: q <= 32'b10111110101010111000001110100001 ;
        130: q <= 32'b10111101000011110001000100101111 ;
        131: q <= 32'b10111111010011001111010101110101 ;
        132: q <= 32'b00111110101011101001101011110000 ;
        133: q <= 32'b00111110101111111110101100101010 ;
        134: q <= 32'b10111110011011101111011011101000 ;
        135: q <= 32'b10111110101111011000011000101010 ;
        136: q <= 32'b10111101101110001101110111011100 ;
        137: q <= 32'b00111110100001101110110100111100 ;
        138: q <= 32'b00111110100100000111110010101100 ;
        139: q <= 32'b10111110011001011000100110111000 ;
        140: q <= 32'b10111110010001111000010000101110 ;
        141: q <= 32'b10111110100100000110101010010000 ;
        142: q <= 32'b00111110101100101101010101111001 ;
        143: q <= 32'b00111110011011011010010010110011 ;
        144: q <= 32'b10111110100010000110100001000100 ;
        145: q <= 32'b00111111001011010010000011110111 ;
        146: q <= 32'b10111111000110101001011100100100 ;
        147: q <= 32'b00111110001101111011010001110111 ;
        148: q <= 32'b10111111010111101011011110011111 ;
        149: q <= 32'b00111110101011101101101001101011 ;
        150: q <= 32'b10111110001000100011100010000011 ;
        151: q <= 32'b00111110100101011100010010000011 ;
        152: q <= 32'b10111110010000011000111110101010 ;
        153: q <= 32'b10111101101111010110110011110100 ;
        154: q <= 32'b00111111001001100010000111101111 ;
        155: q <= 32'b00111110101001101000000111000101 ;
        156: q <= 32'b00111110100111101100011000011110 ;
        157: q <= 32'b10111110010100100011001110100000 ;
        158: q <= 32'b00111110010011001100110111000111 ;
        159: q <= 32'b10111101111111000111100101010111 ;
        160: q <= 32'b00111110001010111110000111110110 ;
        161: q <= 32'b10111110010111100010100100000111 ;
        162: q <= 32'b10111101001000000010001011110010 ;
        163: q <= 32'b10111110001010010101000010111010 ;
        164: q <= 32'b00111110011011010111101100101011 ;
        165: q <= 32'b00111111010100111010101101001111 ;
        166: q <= 32'b10111101101111100011000100000001 ;
        167: q <= 32'b10111110100010111011110111000111 ;
        168: q <= 32'b10111110011010011100000100011101 ;
        169: q <= 32'b10111101011100100100011001011101 ;
        170: q <= 32'b00111110101100001001010000111000 ;
        171: q <= 32'b00111111001010010100011010010011 ;
        172: q <= 32'b00111111000010011011010100001101 ;
        173: q <= 32'b10111101100000000111011110011010 ;
        174: q <= 32'b10111111010101110000111001110100 ;
        175: q <= 32'b00111110100011100000001100110101 ;
        176: q <= 32'b00111100000100100010101011111010 ;
        177: q <= 32'b00111110110100111010110011000111 ;
        178: q <= 32'b10111110100111001011110100000101 ;
        179: q <= 32'b00111110001101110111110101101000 ;
        180: q <= 32'b10111110010101101111010011000100 ;
        181: q <= 32'b00111100010011110101100011101000 ;
        182: q <= 32'b00111110110101000010010101110010 ;
        183: q <= 32'b10111110000100100111010001001111 ;
        184: q <= 32'b10111110010011101001110100001101 ;
        185: q <= 32'b10111110101010000110000000101111 ;
        186: q <= 32'b10111110010000001011111111100110 ;
        187: q <= 32'b10111110000100110111011011000100 ;
        188: q <= 32'b00000000000000000000000000000000 ;
        189: q <= 32'b00000000000000000000000000000000 ;
        190: q <= 32'b00000000000000000000000000000000 ;
        191: q <= 32'b00000000000000000000000000000000 ;
        192: q <= 32'b00111110100110111111011101100111 ;
        193: q <= 32'b00111110100011110000111111011100 ;
        194: q <= 32'b10111110000001111000100000010011 ;
        195: q <= 32'b00111111001000110100001011011010 ;
        196: q <= 32'b10111011110010000100001011000111 ;
        197: q <= 32'b00111110001101011101111001010001 ;
        198: q <= 32'b10111110101001011000101010100010 ;
        199: q <= 32'b10111110100111000011110111000111 ;
        200: q <= 32'b00111110010011110101100101101010 ;
        201: q <= 32'b10111100011101101101011111110000 ;
        202: q <= 32'b10111111010000001000110001000100 ;
        203: q <= 32'b10111100001011100110000101110010 ;
        204: q <= 32'b00111101101111100000001001110111 ;
        205: q <= 32'b10111110100011101000010110101011 ;
        206: q <= 32'b10111101000000110111000111001001 ;
        207: q <= 32'b00111101100001110001001011011110 ;
        208: q <= 32'b00111101011101010110010010111100 ;
        209: q <= 32'b00111111000110100100001000111101 ;
        210: q <= 32'b00111110100100000111001111101110 ;
        211: q <= 32'b00111101110011010101101000001100 ;
        212: q <= 32'b00111110010101001010100001000010 ;
        213: q <= 32'b00111101010000001001110010100100 ;
        214: q <= 32'b10111110001010101111001110110110 ;
        215: q <= 32'b00111110100010001100000110110101 ;
        216: q <= 32'b10111100100111011001101011000111 ;
        217: q <= 32'b10111101011110110000011001100001 ;
        218: q <= 32'b00111111010101011110111101010111 ;
        219: q <= 32'b00111110000111100101110110000100 ;
        220: q <= 32'b00111110011110111001110001110000 ;
        221: q <= 32'b10111110011100110110111010101000 ;
        222: q <= 32'b00111110000111110111100001110001 ;
        223: q <= 32'b10111111001101000010001001001111 ;
        224: q <= 32'b00111101000101001100110111100101 ;
        225: q <= 32'b10111110100000011001101001000011 ;
        226: q <= 32'b10111100001011000000000011011010 ;
        227: q <= 32'b10111110100110100011101001001001 ;
        228: q <= 32'b00111110101001001110101010011101 ;
        229: q <= 32'b00111110011100111100100110011010 ;
        230: q <= 32'b00111100011101100111001010111101 ;
        231: q <= 32'b00111111000000001001100001111101 ;
        232: q <= 32'b10111110101011100100010101100001 ;
        233: q <= 32'b10111101010110011110100111001010 ;
        234: q <= 32'b00111110100110000111111101101101 ;
        235: q <= 32'b00111111000100101110110011110001 ;
        236: q <= 32'b00111101101110100111110010010001 ;
        237: q <= 32'b10111101111101010110000000001110 ;
        238: q <= 32'b00111110000010011000101111000010 ;
        239: q <= 32'b10111101100010110100100100111110 ;
        240: q <= 32'b10111111000001000001101010010000 ;
        241: q <= 32'b00111110110100001110101000000010 ;
        242: q <= 32'b10111110101111010000100011100010 ;
        243: q <= 32'b00111110001001111011110001111110 ;
        244: q <= 32'b10111101111110111101000000101000 ;
        245: q <= 32'b10111101000111111110101110101000 ;
        246: q <= 32'b10111110101011110110101111001100 ;
        247: q <= 32'b00111111011101100100111100101111 ;
        248: q <= 32'b00111111001001000011110101011100 ;
        249: q <= 32'b10111110011111111010010100000000 ;
        250: q <= 32'b10111110010100100100010010101110 ;
        251: q <= 32'b10111110100101111101110001011101 ;
        252: q <= 32'b00000000000000000000000000000000 ;
        253: q <= 32'b00000000000000000000000000000000 ;
        254: q <= 32'b00000000000000000000000000000000 ;
        255: q <= 32'b00000000000000000000000000000000 ;
        256: q <= 32'b00111110000110001011011100101101 ;
        257: q <= 32'b00111101111011011111000001010111 ;
        258: q <= 32'b10111110010101000100101000011100 ;
        259: q <= 32'b10111101010010110111111100101110 ;
        260: q <= 32'b00111110011001010111011011110111 ;
        261: q <= 32'b00111110101110000010111111110100 ;
        262: q <= 32'b10111110011100010111101110101100 ;
        263: q <= 32'b10111110001011100111100110010101 ;
        264: q <= 32'b00111101011101111101011010111101 ;
        265: q <= 32'b00111110001011101100001010110001 ;
        266: q <= 32'b10111101110110010101011001110100 ;
        267: q <= 32'b10111111001111001111111000110101 ;
        268: q <= 32'b00111101110011101010111010010111 ;
        269: q <= 32'b10111110011101001010000010101011 ;
        270: q <= 32'b00111110111011101000110011010101 ;
        271: q <= 32'b00111110110011011000110111111011 ;
        272: q <= 32'b10111110011100000110100101010111 ;
        273: q <= 32'b10111110000100110100001110111110 ;
        274: q <= 32'b10111111000001101110100000101100 ;
        275: q <= 32'b00111111010101000010001001011011 ;
        276: q <= 32'b00111101111110010000000110111100 ;
        277: q <= 32'b10111101101110000111111101000010 ;
        278: q <= 32'b10111110011010000111110101000010 ;
        279: q <= 32'b00111101111000010011100000000110 ;
        280: q <= 32'b10111101011010010110111110000100 ;
        281: q <= 32'b10111111001011100011001010101111 ;
        282: q <= 32'b00111110110111100101001111010110 ;
        283: q <= 32'b00111110001101111110001101111011 ;
        284: q <= 32'b00111110001010110101001110111101 ;
        285: q <= 32'b10111110000000001010100011011100 ;
        286: q <= 32'b00111110011010101001001111010111 ;
        287: q <= 32'b10111011101110001110101111001011 ;
        288: q <= 32'b00111110111110011010101100010010 ;
        289: q <= 32'b10111110000110001001111010011001 ;
        290: q <= 32'b00111110101011111111001100101010 ;
        291: q <= 32'b00111110010101011111001101000100 ;
        292: q <= 32'b00111110100100000010011100000110 ;
        293: q <= 32'b00111100011101011100101100001111 ;
        294: q <= 32'b00111011101111001110111110010000 ;
        295: q <= 32'b10111110100011111011010010100110 ;
        296: q <= 32'b10111101111101000110110011110011 ;
        297: q <= 32'b10111110111100110010000110101101 ;
        298: q <= 32'b00111110001010101000000001000010 ;
        299: q <= 32'b00111110000100111011011111001001 ;
        300: q <= 32'b10111111000111100011011001111111 ;
        301: q <= 32'b10111101010101100110001000011000 ;
        302: q <= 32'b00111101011110110001011100110100 ;
        303: q <= 32'b00111110000110001101110011000100 ;
        304: q <= 32'b10111110101011010110000011110111 ;
        305: q <= 32'b10111101010110000011001000010010 ;
        306: q <= 32'b10111110011111000101000101011000 ;
        307: q <= 32'b00111101110101000011000011010111 ;
        308: q <= 32'b00111101011000011000011110001010 ;
        309: q <= 32'b00111111000010110001011111110000 ;
        310: q <= 32'b00111110011111001000000011100000 ;
        311: q <= 32'b10111101000011000101101110010000 ;
        312: q <= 32'b10111101010101111110001111011001 ;
        313: q <= 32'b10111101111110001111101110100110 ;
        314: q <= 32'b10111110110111010110100010001010 ;
        315: q <= 32'b10111101110100101000011100000001 ;
        316: q <= 32'b00000000000000000000000000000000 ;
        317: q <= 32'b00000000000000000000000000000000 ;
        318: q <= 32'b00000000000000000000000000000000 ;
        319: q <= 32'b00000000000000000000000000000000 ;
        320: q <= 32'b00111110100000100000100000011111 ;
        321: q <= 32'b10111111001010001001001100100001 ;
        322: q <= 32'b10111101110000011101111000111010 ;
        323: q <= 32'b10111111010000100010011111010100 ;
        324: q <= 32'b00111110011001111110010101010101 ;
        325: q <= 32'b00111110101011100000010111010110 ;
        326: q <= 32'b10111110000111101111011001011011 ;
        327: q <= 32'b10111110101100101001100001111101 ;
        328: q <= 32'b00111101101000001110111100111010 ;
        329: q <= 32'b10111110110101111100000111101110 ;
        330: q <= 32'b10111111011001000001001110100111 ;
        331: q <= 32'b10111110000111101101110101110010 ;
        332: q <= 32'b00111110001100001111110110101110 ;
        333: q <= 32'b10111110001010110110101011100011 ;
        334: q <= 32'b00111101101110001100010111000100 ;
        335: q <= 32'b00111101010100100001111001000001 ;
        336: q <= 32'b10111011110111011010001001000001 ;
        337: q <= 32'b10111110110101111001001101101100 ;
        338: q <= 32'b00111110111100100110101010100011 ;
        339: q <= 32'b00111110000101011000111010101000 ;
        340: q <= 32'b10111110000111000101010100110100 ;
        341: q <= 32'b00111101111010001001001100010000 ;
        342: q <= 32'b10111100111011001100010001001111 ;
        343: q <= 32'b00111110010110001001100000111110 ;
        344: q <= 32'b10111110010011111110011111001101 ;
        345: q <= 32'b10111100011010010101011001110101 ;
        346: q <= 32'b00111110110111110111010101001000 ;
        347: q <= 32'b00111110001010000100100101010100 ;
        348: q <= 32'b00111110101001010000010110010111 ;
        349: q <= 32'b10111110000000000110011010010111 ;
        350: q <= 32'b00111101101001011100100011010000 ;
        351: q <= 32'b00111110101100100010101101011010 ;
        352: q <= 32'b00111101010110100010100011111000 ;
        353: q <= 32'b10111110011100011010000011111111 ;
        354: q <= 32'b10111110001001011110010010011101 ;
        355: q <= 32'b10111110010011001001000110001110 ;
        356: q <= 32'b00111110101011010001110011101111 ;
        357: q <= 32'b10111101000010001101101000101101 ;
        358: q <= 32'b10111110100101010011010011011110 ;
        359: q <= 32'b00111111001100100101110000110001 ;
        360: q <= 32'b10111110000011100110110001110000 ;
        361: q <= 32'b10111100101000011001110110101000 ;
        362: q <= 32'b00111110010000110010000001011001 ;
        363: q <= 32'b10111101111111001011001110000101 ;
        364: q <= 32'b00111101101101010000111100101101 ;
        365: q <= 32'b10111100011101100110000111000001 ;
        366: q <= 32'b10111111010101101010111101111111 ;
        367: q <= 32'b00111110000010110011110011001101 ;
        368: q <= 32'b10111111010101100001011111000111 ;
        369: q <= 32'b00111110111010000111111100100001 ;
        370: q <= 32'b10111110101000011000011110110101 ;
        371: q <= 32'b10111101101101110000111010100111 ;
        372: q <= 32'b00111111011111111101111010000101 ;
        373: q <= 32'b00111110001110011101001011000001 ;
        374: q <= 32'b10111110111000111110011011001011 ;
        375: q <= 32'b00111011111110000001010001110001 ;
        376: q <= 32'b10111110010000100101000111100100 ;
        377: q <= 32'b10111110000101001010001100110011 ;
        378: q <= 32'b00111110110111010000100110100000 ;
        379: q <= 32'b10111110001101011101001111101001 ;
        380: q <= 32'b00000000000000000000000000000000 ;
        381: q <= 32'b00000000000000000000000000000000 ;
        382: q <= 32'b00000000000000000000000000000000 ;
        383: q <= 32'b00000000000000000000000000000000 ;
        384: q <= 32'b00111110011110111001001111000011 ;
        385: q <= 32'b10111111000000100111001101011000 ;
        386: q <= 32'b10111110100001001110101000101111 ;
        387: q <= 32'b00111110000000010101100000111100 ;
        388: q <= 32'b00111110101111000010111001001110 ;
        389: q <= 32'b10111111000100000011000010111100 ;
        390: q <= 32'b10111110011100011111101110101111 ;
        391: q <= 32'b10111110010000101000110001001010 ;
        392: q <= 32'b10111111001101010100101011010101 ;
        393: q <= 32'b10111101111011100110010010001011 ;
        394: q <= 32'b00111101101010010010110100111000 ;
        395: q <= 32'b00111101110110000110010100110110 ;
        396: q <= 32'b00111110100110001011010000011010 ;
        397: q <= 32'b10111110100101110101111101111001 ;
        398: q <= 32'b10111110110110011101011101111101 ;
        399: q <= 32'b00111101101111010000011011000111 ;
        400: q <= 32'b00111101100011111010001101001101 ;
        401: q <= 32'b00111110101001010100000100011100 ;
        402: q <= 32'b10111110101011000101010100011000 ;
        403: q <= 32'b10111110001100010110000010110110 ;
        404: q <= 32'b00111100001100011100100100100011 ;
        405: q <= 32'b00111110001000110010110100001111 ;
        406: q <= 32'b10111110011000010000101110100110 ;
        407: q <= 32'b10111100100101110001011110001110 ;
        408: q <= 32'b10111111011010000011000110001001 ;
        409: q <= 32'b10111110010101000010101111010011 ;
        410: q <= 32'b10111110100110101100100011101010 ;
        411: q <= 32'b00111110100101010110100110100001 ;
        412: q <= 32'b00111101100101101100001111010000 ;
        413: q <= 32'b10111110100100101110001000111101 ;
        414: q <= 32'b00111110001101000111000011001100 ;
        415: q <= 32'b10111100111011010101010110001001 ;
        416: q <= 32'b10111101000000101001111010000001 ;
        417: q <= 32'b10111110000111000111001000110111 ;
        418: q <= 32'b10111100100011110000000001001111 ;
        419: q <= 32'b10111110111000100001001001011100 ;
        420: q <= 32'b00111110000101011010110111101101 ;
        421: q <= 32'b10111110000000000010010010111001 ;
        422: q <= 32'b00111101101011011100011011001010 ;
        423: q <= 32'b10111111000000101011011010111010 ;
        424: q <= 32'b10111110100111011000010010111011 ;
        425: q <= 32'b00111110000110110011000001100101 ;
        426: q <= 32'b00111110100101100101111001010010 ;
        427: q <= 32'b00111111000001010100110000010101 ;
        428: q <= 32'b10111111000101101010011111011001 ;
        429: q <= 32'b10111111001100111101010011100000 ;
        430: q <= 32'b10111101101111110000000000001010 ;
        431: q <= 32'b10111101000111111100001111010011 ;
        432: q <= 32'b10111100011010100011001001101100 ;
        433: q <= 32'b00111110000011100010001111001010 ;
        434: q <= 32'b10111110000011110111111100000100 ;
        435: q <= 32'b00111101111000111000101110111110 ;
        436: q <= 32'b00111111000111000110000001101000 ;
        437: q <= 32'b00111101100010011010001000001110 ;
        438: q <= 32'b10111110101001100000101100000000 ;
        439: q <= 32'b00111101111001010100111100010010 ;
        440: q <= 32'b10111101100100110000011100011110 ;
        441: q <= 32'b10111110001011000001010101111011 ;
        442: q <= 32'b00111110111011000011110000101110 ;
        443: q <= 32'b10111110011001110010100000111110 ;
        444: q <= 32'b00000000000000000000000000000000 ;
        445: q <= 32'b00000000000000000000000000000000 ;
        446: q <= 32'b00000000000000000000000000000000 ;
        447: q <= 32'b00000000000000000000000000000000 ;
        448: q <= 32'b00111110100000111100001001100001 ;
        449: q <= 32'b10111110110011100110011110000011 ;
        450: q <= 32'b10111101001111011001011101010001 ;
        451: q <= 32'b10111111001001001011011001011100 ;
        452: q <= 32'b00111110100000110110111001111011 ;
        453: q <= 32'b00111101111100001110011100110011 ;
        454: q <= 32'b10111101010001010001100000101111 ;
        455: q <= 32'b10111110100001100100100010111000 ;
        456: q <= 32'b10111111010000010111101011011111 ;
        457: q <= 32'b10111101001101111101101000010101 ;
        458: q <= 32'b00111110010100010011001111010101 ;
        459: q <= 32'b10111101110011011110011101110111 ;
        460: q <= 32'b00111101110011000010100111100100 ;
        461: q <= 32'b10111110100100010001111010001110 ;
        462: q <= 32'b00111101111100101100110010101101 ;
        463: q <= 32'b00111110000001110001110001010100 ;
        464: q <= 32'b10111110010111001011100010010001 ;
        465: q <= 32'b10111110101001000000011110011101 ;
        466: q <= 32'b00111110111001000001101000101000 ;
        467: q <= 32'b00111100110001110000001001101100 ;
        468: q <= 32'b00111101111010110101111100111111 ;
        469: q <= 32'b10111111001101111000100010011110 ;
        470: q <= 32'b10111101110101000001100000101101 ;
        471: q <= 32'b00111110000000001101011110001110 ;
        472: q <= 32'b00111101011011000011111001001100 ;
        473: q <= 32'b00111100101101110000001100001101 ;
        474: q <= 32'b10111110100100000100111011001100 ;
        475: q <= 32'b00111110101001001110001110000000 ;
        476: q <= 32'b00111110001111110111001011100001 ;
        477: q <= 32'b10111110011010000101011010000111 ;
        478: q <= 32'b00111101100100111010001000100011 ;
        479: q <= 32'b10111100111001010110011010111000 ;
        480: q <= 32'b00111010100000010010001101011100 ;
        481: q <= 32'b10111110000100000110110011001110 ;
        482: q <= 32'b00111111010010110000101101111110 ;
        483: q <= 32'b00111110000110111101011100111010 ;
        484: q <= 32'b00111110010000100101001010000010 ;
        485: q <= 32'b10111101011010101011000001001110 ;
        486: q <= 32'b10111100010001010011111010100111 ;
        487: q <= 32'b00111110111110110110001001111011 ;
        488: q <= 32'b10111110101000011111101111111010 ;
        489: q <= 32'b10111101001101111101010000001110 ;
        490: q <= 32'b00111110100111111000101110110010 ;
        491: q <= 32'b10111110010011100100010000100010 ;
        492: q <= 32'b10111110110110101010010001100010 ;
        493: q <= 32'b00111101000010110110010011111011 ;
        494: q <= 32'b10111111001000000110001101101100 ;
        495: q <= 32'b00111100011110100111101010110001 ;
        496: q <= 32'b00111110011111011100111100001001 ;
        497: q <= 32'b10111110111100111100011111001100 ;
        498: q <= 32'b10111101110110010010011010100101 ;
        499: q <= 32'b00111111010110000010111000001000 ;
        500: q <= 32'b10111101100100000000011111101011 ;
        501: q <= 32'b00111011001100001111011001011111 ;
        502: q <= 32'b00111110001010001010001111101000 ;
        503: q <= 32'b10111100010101011001001110010011 ;
        504: q <= 32'b10111110000011001011100011101000 ;
        505: q <= 32'b10111101110100011001111101101001 ;
        506: q <= 32'b10111100101100101101100100001111 ;
        507: q <= 32'b10111101100111111011101100111001 ;
        508: q <= 32'b00000000000000000000000000000000 ;
        509: q <= 32'b00000000000000000000000000000000 ;
        510: q <= 32'b00000000000000000000000000000000 ;
        511: q <= 32'b00000000000000000000000000000000 ;
        512: q <= 32'b00111110101011101010111100100101 ;
        513: q <= 32'b00111111000011101010001101010001 ;
        514: q <= 32'b10111101101110010101101101011100 ;
        515: q <= 32'b10111111011011100100001110010011 ;
        516: q <= 32'b10111100110001100100101010101110 ;
        517: q <= 32'b00111110101101111101101011111000 ;
        518: q <= 32'b10111110100000011001100011110100 ;
        519: q <= 32'b10111110101111100010000111000110 ;
        520: q <= 32'b00111110000111111110111000100000 ;
        521: q <= 32'b10111110010000000011001111010011 ;
        522: q <= 32'b10111111010100011000000100011100 ;
        523: q <= 32'b10111110101010100001010011101000 ;
        524: q <= 32'b00111110011011111101000000101100 ;
        525: q <= 32'b10111110000111000110001000110111 ;
        526: q <= 32'b10111101000011111111111001010010 ;
        527: q <= 32'b00111100010000000101111000010100 ;
        528: q <= 32'b10111110011100010000111111101011 ;
        529: q <= 32'b00111111000100101101000001110010 ;
        530: q <= 32'b00111110111111010101101100011010 ;
        531: q <= 32'b00111101111111000011100010110111 ;
        532: q <= 32'b10111100101101110111010000100000 ;
        533: q <= 32'b00111101010001100101101010111011 ;
        534: q <= 32'b00111101010001110100111011101010 ;
        535: q <= 32'b00111110100011100000000010000101 ;
        536: q <= 32'b10111110000101110001010011110010 ;
        537: q <= 32'b00111100110111000101101001010110 ;
        538: q <= 32'b10111111010010100110110110010100 ;
        539: q <= 32'b00111110101110010101111000110110 ;
        540: q <= 32'b00111110011110100111000101000110 ;
        541: q <= 32'b10111110101111101100000000001001 ;
        542: q <= 32'b00111110011001000010010110000001 ;
        543: q <= 32'b10111111001011001100000110111011 ;
        544: q <= 32'b00111011111111101110101010010001 ;
        545: q <= 32'b10111110100111111010001100010101 ;
        546: q <= 32'b00111100110100000011011011001100 ;
        547: q <= 32'b10111110100101111001110101110100 ;
        548: q <= 32'b00111110100011100010000111001000 ;
        549: q <= 32'b10111101001001111110001010010101 ;
        550: q <= 32'b00111101000001000000011111100010 ;
        551: q <= 32'b10111111000101010101001010000101 ;
        552: q <= 32'b10111110010100101001101000101111 ;
        553: q <= 32'b10111110000110111100110101111010 ;
        554: q <= 32'b00111110100101101111010101010101 ;
        555: q <= 32'b10111110111100010000010100001011 ;
        556: q <= 32'b00111110001011110000000101111101 ;
        557: q <= 32'b10111101110011011011010101101011 ;
        558: q <= 32'b00111101101010001011000000010101 ;
        559: q <= 32'b10111101000110010010111110000011 ;
        560: q <= 32'b10111111000110001011001101011000 ;
        561: q <= 32'b10111111011101011010100110101011 ;
        562: q <= 32'b10111110110001110000101101000101 ;
        563: q <= 32'b10111110000001001010101101001101 ;
        564: q <= 32'b10111110010100001101111001001101 ;
        565: q <= 32'b10111101010001110010111010001101 ;
        566: q <= 32'b10111110111111010001110011111110 ;
        567: q <= 32'b10111110100100010000001001000000 ;
        568: q <= 32'b10111111000001000001000001101111 ;
        569: q <= 32'b10111110100011000000110001101001 ;
        570: q <= 32'b10111110100101010101010110010101 ;
        571: q <= 32'b10111110101101010000111010011111 ;
        572: q <= 32'b00000000000000000000000000000000 ;
        573: q <= 32'b00000000000000000000000000000000 ;
        574: q <= 32'b00000000000000000000000000000000 ;
        575: q <= 32'b00000000000000000000000000000000 ;
        576: q <= 32'b00111110001110001101111001001001 ;
        577: q <= 32'b00111110101101001001011100110010 ;
        578: q <= 32'b10111110010101010011000110100001 ;
        579: q <= 32'b10111100110101111011110010100000 ;
        580: q <= 32'b00111101100001011001101111101011 ;
        581: q <= 32'b10111110101110000011100100001001 ;
        582: q <= 32'b10111110001001111011011000110011 ;
        583: q <= 32'b10111101110111000001100101010010 ;
        584: q <= 32'b10111101000100101000000101000100 ;
        585: q <= 32'b10111111010000001011100110101011 ;
        586: q <= 32'b00111110001100101001101111010101 ;
        587: q <= 32'b00111011110011111011010011000001 ;
        588: q <= 32'b10111110010011101001010101000100 ;
        589: q <= 32'b10111110000010101101010000100010 ;
        590: q <= 32'b00111110100010100100111000001000 ;
        591: q <= 32'b10111100001100000100110100111011 ;
        592: q <= 32'b00111100101010010001100000010111 ;
        593: q <= 32'b10111110001101110010111110110100 ;
        594: q <= 32'b00111110000111111011011100000101 ;
        595: q <= 32'b00111110000101111101000010010100 ;
        596: q <= 32'b10111110110001100111010111000101 ;
        597: q <= 32'b10111101111001101110100010111011 ;
        598: q <= 32'b00111110101001100001001110011111 ;
        599: q <= 32'b00111110001000001110011011010010 ;
        600: q <= 32'b10111101001011011101000111001000 ;
        601: q <= 32'b10111110010000110100001011001111 ;
        602: q <= 32'b00111110101010001110100101100001 ;
        603: q <= 32'b00111110100111100111010101001110 ;
        604: q <= 32'b00111110000100001001111100001001 ;
        605: q <= 32'b10111110100100111110111100010110 ;
        606: q <= 32'b00111111011110000000100000010110 ;
        607: q <= 32'b10111111010011010000110010000001 ;
        608: q <= 32'b10111010001111000101011011110101 ;
        609: q <= 32'b10111101111001010110011110101011 ;
        610: q <= 32'b00111101101101110110011111010110 ;
        611: q <= 32'b10111110001100011100011000011100 ;
        612: q <= 32'b00111110011110100010100011000011 ;
        613: q <= 32'b10111110010110101001101100101110 ;
        614: q <= 32'b10111110010010010000111001100110 ;
        615: q <= 32'b10111110100011010010101110101110 ;
        616: q <= 32'b10111110100011100101111101111111 ;
        617: q <= 32'b00111101001001100111110001110110 ;
        618: q <= 32'b00111110011001011001000101110110 ;
        619: q <= 32'b00111101101001110011101111000010 ;
        620: q <= 32'b00111101001001010011010011111001 ;
        621: q <= 32'b10111110000011000000100001101111 ;
        622: q <= 32'b10111111000000000001011110100101 ;
        623: q <= 32'b10111111000011000001000100110100 ;
        624: q <= 32'b00111110010101010000111011000111 ;
        625: q <= 32'b00111110001001100011011010011100 ;
        626: q <= 32'b10111110011001111111011011000100 ;
        627: q <= 32'b00111011101111110101101000111100 ;
        628: q <= 32'b00111111001100001011011001111101 ;
        629: q <= 32'b00111100001010011011010010100101 ;
        630: q <= 32'b00111110011010101100000100011011 ;
        631: q <= 32'b00111110000100110001110000100110 ;
        632: q <= 32'b00111110000100101101100011100110 ;
        633: q <= 32'b10111110001111000100111110100000 ;
        634: q <= 32'b10111110101100110100011010011111 ;
        635: q <= 32'b10111110011111110111001010010001 ;
        636: q <= 32'b00000000000000000000000000000000 ;
        637: q <= 32'b00000000000000000000000000000000 ;
        638: q <= 32'b00000000000000000000000000000000 ;
        639: q <= 32'b00000000000000000000000000000000 ;
        640: q <= 32'b00111110101110010101110000010001 ;
        641: q <= 32'b10111111000011000001000000001001 ;
        642: q <= 32'b00111101001001110100000101100011 ;
        643: q <= 32'b10111111000001111101000101001001 ;
        644: q <= 32'b00111110010101001111111001101010 ;
        645: q <= 32'b10111111010010100100111011010110 ;
        646: q <= 32'b10111110110001001000001001001011 ;
        647: q <= 32'b10111110101001000010011101000111 ;
        648: q <= 32'b10111101000000111100000101111110 ;
        649: q <= 32'b10111110000000001011101110110110 ;
        650: q <= 32'b00111110100111000110010110001010 ;
        651: q <= 32'b10111110010010101110101000010111 ;
        652: q <= 32'b00111101000011010001011010111111 ;
        653: q <= 32'b10111110100000001001100000100000 ;
        654: q <= 32'b00111110101010001010101111001011 ;
        655: q <= 32'b00111101000001110001001001011101 ;
        656: q <= 32'b10111110111111011100110011110001 ;
        657: q <= 32'b10111111000110100110010110011111 ;
        658: q <= 32'b10111111001100011011100100100011 ;
        659: q <= 32'b00111110001011001111001000010100 ;
        660: q <= 32'b00111110011000010100110010101111 ;
        661: q <= 32'b00111110010110011010000001100100 ;
        662: q <= 32'b10111110000101100111000000100101 ;
        663: q <= 32'b00111110001011011001111100010000 ;
        664: q <= 32'b10111101100110101010011001001001 ;
        665: q <= 32'b10111100100001110110111001100010 ;
        666: q <= 32'b00111111001100110011010011111000 ;
        667: q <= 32'b00111110101010100011111110101001 ;
        668: q <= 32'b00111110101001000011011100001110 ;
        669: q <= 32'b10111110100011000111010000101000 ;
        670: q <= 32'b00111110001100110111000011000011 ;
        671: q <= 32'b00111101010110001011001000110000 ;
        672: q <= 32'b10111101100100111111010010111100 ;
        673: q <= 32'b10111101110000111101011001100001 ;
        674: q <= 32'b10111101111011111111111100100010 ;
        675: q <= 32'b10111110101000110010100110011001 ;
        676: q <= 32'b00111110101100111111010001110100 ;
        677: q <= 32'b10111110101110001111110101010001 ;
        678: q <= 32'b10111110101001000011110010101101 ;
        679: q <= 32'b10111110101001111011101011101001 ;
        680: q <= 32'b10111110101111000001100001001110 ;
        681: q <= 32'b00111101111011000011000010010000 ;
        682: q <= 32'b00111110100011001001110011011100 ;
        683: q <= 32'b10111110101010010101001010001011 ;
        684: q <= 32'b00111111000010000101111111011010 ;
        685: q <= 32'b10111110010011000101111000011011 ;
        686: q <= 32'b00111110110111100101110100011110 ;
        687: q <= 32'b10111101100001000000111001100000 ;
        688: q <= 32'b10111111001011110110100111111010 ;
        689: q <= 32'b10111111001110110010000111110000 ;
        690: q <= 32'b10111110100100101000101111101111 ;
        691: q <= 32'b00111101010101101010101110110001 ;
        692: q <= 32'b10111110100001101110111001111001 ;
        693: q <= 32'b10111100011110110101110101101001 ;
        694: q <= 32'b10111110100001000011111000000010 ;
        695: q <= 32'b00111110010001101100010000100101 ;
        696: q <= 32'b00111111010001011011001111001010 ;
        697: q <= 32'b10111110000110100010111100110101 ;
        698: q <= 32'b00111110001000000111100001011101 ;
        699: q <= 32'b10111110110011111000111110010011 ;
        700: q <= 32'b00000000000000000000000000000000 ;
        701: q <= 32'b00000000000000000000000000000000 ;
        702: q <= 32'b00000000000000000000000000000000 ;
        703: q <= 32'b00000000000000000000000000000000 ;
        704: q <= 32'b00111101111110011100110001101011 ;
        705: q <= 32'b10111110010000000111100000100001 ;
        706: q <= 32'b00111101000000101000100011001011 ;
        707: q <= 32'b10111110101110100001100000000110 ;
        708: q <= 32'b00111110001001001010001110101110 ;
        709: q <= 32'b00111110000101110101100110110010 ;
        710: q <= 32'b10111110001100011010111110101000 ;
        711: q <= 32'b10111110101010001110000000000101 ;
        712: q <= 32'b00111110101001100010011011110111 ;
        713: q <= 32'b10111110100001101011110010111010 ;
        714: q <= 32'b00111101100000011001110001110000 ;
        715: q <= 32'b10111110000111111000010110000101 ;
        716: q <= 32'b10111100100010001000011000100101 ;
        717: q <= 32'b10111110000110110010000111010001 ;
        718: q <= 32'b00111101110101000111010011111011 ;
        719: q <= 32'b00111110001010101001010111110011 ;
        720: q <= 32'b10111101100001101000001000111011 ;
        721: q <= 32'b00111111000001110101010101101011 ;
        722: q <= 32'b10111110101100011000010011001010 ;
        723: q <= 32'b10111100100001101110111001001001 ;
        724: q <= 32'b00111110000100110001001110101011 ;
        725: q <= 32'b10111111001111111111111010101101 ;
        726: q <= 32'b00111101010001111000000010011001 ;
        727: q <= 32'b00111101100000000100001101101100 ;
        728: q <= 32'b00111101110000011010010001001100 ;
        729: q <= 32'b10111110001001110000010110111000 ;
        730: q <= 32'b10111111000100011111010100010110 ;
        731: q <= 32'b00111110100000010101010010010011 ;
        732: q <= 32'b00111110100011100101110111001100 ;
        733: q <= 32'b10111110101010010000010011111010 ;
        734: q <= 32'b00111110100010000010010100000010 ;
        735: q <= 32'b10111011010101101111110110111101 ;
        736: q <= 32'b00111110010001001001011000100000 ;
        737: q <= 32'b10111110001100001011110101100000 ;
        738: q <= 32'b10111110000010111100010110100100 ;
        739: q <= 32'b10111101101111001010011101110000 ;
        740: q <= 32'b00111110100100000010010010000101 ;
        741: q <= 32'b00111111010001100011010000011011 ;
        742: q <= 32'b10111110000000110100101101001011 ;
        743: q <= 32'b10111110011111010100111001001000 ;
        744: q <= 32'b10111110010000011100101100100111 ;
        745: q <= 32'b00111100111010011001000110110010 ;
        746: q <= 32'b00111110001101111010000001100110 ;
        747: q <= 32'b00111111000110101011111001110101 ;
        748: q <= 32'b10111111010000000011100000010010 ;
        749: q <= 32'b10111011110011100001001101000111 ;
        750: q <= 32'b00111110101110000011101100111110 ;
        751: q <= 32'b10111110000000001100011011000010 ;
        752: q <= 32'b00111110101001101010011110111111 ;
        753: q <= 32'b10111111001011000110110110001001 ;
        754: q <= 32'b10111110100100110100001000111101 ;
        755: q <= 32'b10111110000100001100001000011111 ;
        756: q <= 32'b10111101111000011001100110100010 ;
        757: q <= 32'b00111110010000100110110111101001 ;
        758: q <= 32'b10111110101010001101000100110110 ;
        759: q <= 32'b00111110110100001110010100010100 ;
        760: q <= 32'b00111111010100101111011000011100 ;
        761: q <= 32'b10111110001011111100010001010111 ;
        762: q <= 32'b10111110101110001001101011100011 ;
        763: q <= 32'b10111110011011011000111011010011 ;
        764: q <= 32'b00000000000000000000000000000000 ;
        765: q <= 32'b00000000000000000000000000000000 ;
        766: q <= 32'b00000000000000000000000000000000 ;
        767: q <= 32'b00000000000000000000000000000000 ;
        768: q <= 32'b00111101101100100111000001011001 ;
        769: q <= 32'b00111110011101000000101001010101 ;
        770: q <= 32'b10111101011001111110010100011101 ;
        771: q <= 32'b10111110001000000111010100110001 ;
        772: q <= 32'b10111101010010100100100101010011 ;
        773: q <= 32'b10111111000000001101111110111101 ;
        774: q <= 32'b10111110000001100011001101101110 ;
        775: q <= 32'b10111101111010000001111101001010 ;
        776: q <= 32'b10111110110111101101111110010011 ;
        777: q <= 32'b10111101010001011011101010100011 ;
        778: q <= 32'b10111101100011011010100111011101 ;
        779: q <= 32'b10111110000110010110011000000010 ;
        780: q <= 32'b10111101001111001001110011000010 ;
        781: q <= 32'b10111110100010100010001011101000 ;
        782: q <= 32'b10111110011110100000100110110100 ;
        783: q <= 32'b10111100110010100101101001010100 ;
        784: q <= 32'b10111110010011000100111101111110 ;
        785: q <= 32'b10111110011101110100011001010100 ;
        786: q <= 32'b10111110110100001010100011010101 ;
        787: q <= 32'b00111100100111100011111101010000 ;
        788: q <= 32'b00111101001111010111010010100011 ;
        789: q <= 32'b10111110001000110010011101111000 ;
        790: q <= 32'b00111111001100011110011010010010 ;
        791: q <= 32'b00111111011110111011111101100100 ;
        792: q <= 32'b00111100100110100001111000100011 ;
        793: q <= 32'b10111101110101000000110100000100 ;
        794: q <= 32'b10111110111000000010110111110010 ;
        795: q <= 32'b00111101110000010011110101000001 ;
        796: q <= 32'b00111110100111011000011100101000 ;
        797: q <= 32'b10111110100110000001100011011100 ;
        798: q <= 32'b00111110011110011100000101000100 ;
        799: q <= 32'b00111101010011001111000110000001 ;
        800: q <= 32'b10111110000111111110110100010010 ;
        801: q <= 32'b10111111010100100010011000000100 ;
        802: q <= 32'b10111110001000010001010011101110 ;
        803: q <= 32'b00111110111111000101011101001010 ;
        804: q <= 32'b00111110011011101101111100011000 ;
        805: q <= 32'b00111101110000000010110101000000 ;
        806: q <= 32'b00111101010010100010011111011111 ;
        807: q <= 32'b00111110101100011110010101001110 ;
        808: q <= 32'b10111110101010100111110001010101 ;
        809: q <= 32'b10111110111101011101101110010011 ;
        810: q <= 32'b00111101111101101111110000111110 ;
        811: q <= 32'b10111101011001100101010101100100 ;
        812: q <= 32'b10111110110100111110001111001000 ;
        813: q <= 32'b00111100100000101110010111101111 ;
        814: q <= 32'b10111100000111010100110011111110 ;
        815: q <= 32'b00111011111010001011010110111000 ;
        816: q <= 32'b10111111000010001010010111101001 ;
        817: q <= 32'b10111101001111100011101100111110 ;
        818: q <= 32'b10111110100011111001011101000111 ;
        819: q <= 32'b10111101100001110010111110001000 ;
        820: q <= 32'b00111100111000000101101111011110 ;
        821: q <= 32'b10111100100011011000000100011101 ;
        822: q <= 32'b10111110110010111000101100000010 ;
        823: q <= 32'b10111100000000100101111011010101 ;
        824: q <= 32'b00111101101000101000001100010111 ;
        825: q <= 32'b10111110011010101100010011100100 ;
        826: q <= 32'b10111110001111111001100001100110 ;
        827: q <= 32'b10111110000111000001000110000010 ;
        828: q <= 32'b00000000000000000000000000000000 ;
        829: q <= 32'b00000000000000000000000000000000 ;
        830: q <= 32'b00000000000000000000000000000000 ;
        831: q <= 32'b00000000000000000000000000000000 ;
        832: q <= 32'b00111110001010111010111111010101 ;
        833: q <= 32'b00111110110001111011011011111001 ;
        834: q <= 32'b00111111010010001001011001100010 ;
        835: q <= 32'b10111100110110111000011100111011 ;
        836: q <= 32'b00111110000110101100000010000100 ;
        837: q <= 32'b00111110100011101100101001010101 ;
        838: q <= 32'b10111110101100000011110001000011 ;
        839: q <= 32'b10111110101001001110000111011111 ;
        840: q <= 32'b10111110010011011100100000001010 ;
        841: q <= 32'b00111101001001001010001111111100 ;
        842: q <= 32'b00111101100001010001011101101100 ;
        843: q <= 32'b10111100001000111110000101001101 ;
        844: q <= 32'b00111111001011100011001111000000 ;
        845: q <= 32'b10111101111000111001100110110011 ;
        846: q <= 32'b00111110100001000111000011011011 ;
        847: q <= 32'b00111110000010100010111011000100 ;
        848: q <= 32'b10111101101001101001110111101010 ;
        849: q <= 32'b10111110100010000110110111110110 ;
        850: q <= 32'b10111110111001001101000110101100 ;
        851: q <= 32'b00111101100011000110101110010010 ;
        852: q <= 32'b10111111001100101111100111101010 ;
        853: q <= 32'b00111100101100100010001100000101 ;
        854: q <= 32'b00111111000010110010111001110001 ;
        855: q <= 32'b00111101011110001011110101111101 ;
        856: q <= 32'b10111101010110110011011011101101 ;
        857: q <= 32'b00111100010001010100111010110100 ;
        858: q <= 32'b00111110011110001001010010111100 ;
        859: q <= 32'b00111110001110010011111100011010 ;
        860: q <= 32'b00111110001111111011011011100101 ;
        861: q <= 32'b10111110000001100010111101010001 ;
        862: q <= 32'b00111110010011000010000001001011 ;
        863: q <= 32'b00111101000110100000110001101000 ;
        864: q <= 32'b10111101011010110000110110000001 ;
        865: q <= 32'b10111101110100101100001010100010 ;
        866: q <= 32'b10111110101100000001101001100001 ;
        867: q <= 32'b10111110101011111011110100000101 ;
        868: q <= 32'b00111110001101101000101111100111 ;
        869: q <= 32'b10111110001011110010000110000101 ;
        870: q <= 32'b10111101000000001101000101100001 ;
        871: q <= 32'b00111111000010011100111100100001 ;
        872: q <= 32'b10111110100010001110011101010011 ;
        873: q <= 32'b00111101100100100000101000011101 ;
        874: q <= 32'b00111110101000100110000101000000 ;
        875: q <= 32'b10111110000011010100000001100100 ;
        876: q <= 32'b10111111001011011001001000000001 ;
        877: q <= 32'b10111110001111111101101010111011 ;
        878: q <= 32'b10111110011010001010101100101101 ;
        879: q <= 32'b00111101110001010100111000001101 ;
        880: q <= 32'b00111110010110010100101011000110 ;
        881: q <= 32'b10111101101001000001001010001110 ;
        882: q <= 32'b10111110010010110001000010000100 ;
        883: q <= 32'b10111101011011111110001101101011 ;
        884: q <= 32'b10111101100111110110110101111001 ;
        885: q <= 32'b00111110001111110000001000011010 ;
        886: q <= 32'b00111110110100011111000100010110 ;
        887: q <= 32'b00111111011000001010100100001100 ;
        888: q <= 32'b00111110101110110101111010110001 ;
        889: q <= 32'b10111110101000010111101011100000 ;
        890: q <= 32'b10111110010011110011111101011110 ;
        891: q <= 32'b10111110100110111101100101100101 ;
        892: q <= 32'b00000000000000000000000000000000 ;
        893: q <= 32'b00000000000000000000000000000000 ;
        894: q <= 32'b00000000000000000000000000000000 ;
        895: q <= 32'b00000000000000000000000000000000 ;
        896: q <= 32'b00111110010111110011101111001111 ;
        897: q <= 32'b00111110101010010100101101001000 ;
        898: q <= 32'b00111111000101011000010000111111 ;
        899: q <= 32'b00111101111100101110100010000101 ;
        900: q <= 32'b00111110011101001101100001110110 ;
        901: q <= 32'b10111110110010011111010100100011 ;
        902: q <= 32'b10111110100110110011001011000110 ;
        903: q <= 32'b10111110100101010101101100111000 ;
        904: q <= 32'b00111110100000100010100011110000 ;
        905: q <= 32'b00111101111011011110011010011101 ;
        906: q <= 32'b10111111001000010111101011001111 ;
        907: q <= 32'b00111101001010001001111010101001 ;
        908: q <= 32'b00111110001011110111001111100001 ;
        909: q <= 32'b10111110011110100001000100100111 ;
        910: q <= 32'b10111110100111100000000000011101 ;
        911: q <= 32'b10111100101100011011010000000101 ;
        912: q <= 32'b10111110000110111111110101001000 ;
        913: q <= 32'b10111110100100101000001011100001 ;
        914: q <= 32'b10111110110010101010001010100110 ;
        915: q <= 32'b00111011110000100111110001010000 ;
        916: q <= 32'b00111110001010010011010010110001 ;
        917: q <= 32'b10111101111000011011010111000100 ;
        918: q <= 32'b10111110100111011010011111001101 ;
        919: q <= 32'b00111101111010101101111111111100 ;
        920: q <= 32'b00111101001101001101010001101011 ;
        921: q <= 32'b00111101000010001011110110001010 ;
        922: q <= 32'b00111101100110011010000000011110 ;
        923: q <= 32'b00111110010111100001000100001110 ;
        924: q <= 32'b00111110001000010111000011110001 ;
        925: q <= 32'b10111110011010000101110000000100 ;
        926: q <= 32'b10111100100001101010110011111101 ;
        927: q <= 32'b10111110000000011101011010011101 ;
        928: q <= 32'b00111111000101000101110100011101 ;
        929: q <= 32'b10111110010010111100001001001000 ;
        930: q <= 32'b10111110010110010010000000010111 ;
        931: q <= 32'b00111110111011100111001011011010 ;
        932: q <= 32'b00111110100001010110111011100011 ;
        933: q <= 32'b00111110010101011010110101111000 ;
        934: q <= 32'b00111100100010110110110001001111 ;
        935: q <= 32'b10111110011000011100001111111001 ;
        936: q <= 32'b10111110010001001000010000000010 ;
        937: q <= 32'b00111110000001101010110100010111 ;
        938: q <= 32'b00111110000100100011001000111011 ;
        939: q <= 32'b00111101010100000001001000101100 ;
        940: q <= 32'b00111101100001111111100011110001 ;
        941: q <= 32'b10111110000101001001110011010111 ;
        942: q <= 32'b10111111000100000100010000010101 ;
        943: q <= 32'b00111101100111111011010000000000 ;
        944: q <= 32'b00111110010110101011110100011010 ;
        945: q <= 32'b10111111001011110110110100110110 ;
        946: q <= 32'b10111110011101101101001100100000 ;
        947: q <= 32'b00111111000011100100110101100001 ;
        948: q <= 32'b00111111001010111011110100001101 ;
        949: q <= 32'b00111100110000000111000001101000 ;
        950: q <= 32'b10111110101000110101111001110001 ;
        951: q <= 32'b00111110000110111101011110011010 ;
        952: q <= 32'b00111101101110011010101100101101 ;
        953: q <= 32'b10111110100011100110000011001111 ;
        954: q <= 32'b10111110110001011001001010011110 ;
        955: q <= 32'b10111110101001000010111001111010 ;
        956: q <= 32'b00000000000000000000000000000000 ;
        957: q <= 32'b00000000000000000000000000000000 ;
        958: q <= 32'b00000000000000000000000000000000 ;
        959: q <= 32'b00000000000000000000000000000000 ;
        960: q <= 32'b00111110100000011110001000000110 ;
        961: q <= 32'b00111110100100001101100000110111 ;
        962: q <= 32'b00111101101111110010110010011000 ;
        963: q <= 32'b10111110011001100110011111111100 ;
        964: q <= 32'b00111110011001010001001110000110 ;
        965: q <= 32'b10111111000010110010111111011001 ;
        966: q <= 32'b10111110011111101111010100110001 ;
        967: q <= 32'b10111110010110110000001010000000 ;
        968: q <= 32'b00111101100011110001010111111101 ;
        969: q <= 32'b10111111010000111100101011001000 ;
        970: q <= 32'b00111110000011111010101001100110 ;
        971: q <= 32'b00111110101000110111001001001100 ;
        972: q <= 32'b00111101110100001111001110101101 ;
        973: q <= 32'b10111110100110101000101001101000 ;
        974: q <= 32'b10111111000101111101111001110111 ;
        975: q <= 32'b00111111001000111001001011000010 ;
        976: q <= 32'b10111110000001101110000000011010 ;
        977: q <= 32'b10111110011010100101101001011011 ;
        978: q <= 32'b00111110110110101110111010100110 ;
        979: q <= 32'b10111110010111000001111010001110 ;
        980: q <= 32'b00111110010111000110001111001001 ;
        981: q <= 32'b10111110100100010011100001100110 ;
        982: q <= 32'b10111110010111101100010101100010 ;
        983: q <= 32'b00111110010110100001101111100100 ;
        984: q <= 32'b10111110011010011101100110110000 ;
        985: q <= 32'b00111110010011110000010110100101 ;
        986: q <= 32'b10111110101010000000101011111010 ;
        987: q <= 32'b00111110101010000111110011111111 ;
        988: q <= 32'b00111101110111111110111111111001 ;
        989: q <= 32'b10111110100010010001111010000110 ;
        990: q <= 32'b00111110000111100001011000110110 ;
        991: q <= 32'b00111101111011111111111001010000 ;
        992: q <= 32'b00111111000010100100111000000011 ;
        993: q <= 32'b10111110001001100011100110001000 ;
        994: q <= 32'b00111111000001001110000011001100 ;
        995: q <= 32'b00111110010111011001101010100010 ;
        996: q <= 32'b00111110010001010110010000000001 ;
        997: q <= 32'b00111110000101010100100000100111 ;
        998: q <= 32'b00111100100111011111000111001101 ;
        999: q <= 32'b10111101011010001101100011110111 ;
        1000: q <= 32'b10111101110010100100011100001000 ;
        1001: q <= 32'b10111111000100010111101010101100 ;
        1002: q <= 32'b00111110001011001010011011110111 ;
        1003: q <= 32'b00111101100001000000110100101000 ;
        1004: q <= 32'b00111110010101011110100000011110 ;
        1005: q <= 32'b10111101110000000010011010010000 ;
        1006: q <= 32'b00111101101001001001101010100001 ;
        1007: q <= 32'b10111111010001011000000001110111 ;
        1008: q <= 32'b10111111000110100100110001111101 ;
        1009: q <= 32'b10111110010010000111111101001110 ;
        1010: q <= 32'b10111101111010111100011000110111 ;
        1011: q <= 32'b10111101100111000001010000101110 ;
        1012: q <= 32'b10111101110110011100100001010010 ;
        1013: q <= 32'b00111111000001111101000101110110 ;
        1014: q <= 32'b00111101110111101011011101100110 ;
        1015: q <= 32'b00111110000100101101100111011101 ;
        1016: q <= 32'b00111101111111110111001011001101 ;
        1017: q <= 32'b10111110011001010000100110111100 ;
        1018: q <= 32'b00111111000001000011101100000100 ;
        1019: q <= 32'b10111110100000001101111000001110 ;
        1020: q <= 32'b00000000000000000000000000000000 ;
        1021: q <= 32'b00000000000000000000000000000000 ;
        1022: q <= 32'b00000000000000000000000000000000 ;
        1023: q <= 32'b00000000000000000000000000000000 ;
        default: q <= 32'b00000000000000000000000000000000;
    endcase
end

endmodule
